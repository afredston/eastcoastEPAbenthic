
Search Parameters:Biogeographic Province in (Carolinian))	
Data Group	Sampling Year	Station Name	Sampling Collection Date	Latitude Decimal Degrees	Longitude Decimal Degrees	Visit Number	Station Depth	Depth Units	
EMAP Carolinian Province	1994	CP94001	15-AUG-1994	27.201	-80.176	1	1.2	m	
EMAP Carolinian Province	1994	CP94002	15-AUG-1994	27.214	-80.22	1	3.0	m	
EMAP Carolinian Province	1994	CP94003	16-AUG-1994	27.405	-80.288	1	1.7	m	
EMAP Carolinian Province	1994	CP94004	16-AUG-1994	27.535	-80.33	1	1.0	m	
EMAP Carolinian Province	1994	CP94005	02-AUG-1994	27.679	-80.386	1	0.5	m	
EMAP Carolinian Province	1994	CP94006	03-AUG-1994	27.897	-80.503	1	1.4	m	
EMAP Carolinian Province	1994	CP94007	16-AUG-1994	27.917	-80.507	1	1.4	m	
EMAP Carolinian Province	1994	CP94008	03-AUG-1994	27.995	-80.553	1	1.5	m	
EMAP Carolinian Province	1994	CP94009	01-AUG-1994	28.161	-80.619	1	2.7	m	
EMAP Carolinian Province	1994	CP94010	17-AUG-1994	28.257	-80.675	1	4.0	m	
EMAP Carolinian Province	1994	CP94011	17-AUG-1994	28.503	-80.748	1	1.3	m	
EMAP Carolinian Province	1994	CP94012	18-AUG-1994	28.713	-80.794	1	1.5	m	
EMAP Carolinian Province	1994	CP94013	18-AUG-1994	28.722	-80.803	1	1.5	m	
EMAP Carolinian Province	1994	CP94014	18-AUG-1994	28.852	-80.791	1	1.7	m	
EMAP Carolinian Province	1994	CP94016	08-AUG-1994	30.134	-81.626	1	1.5	m	
EMAP Carolinian Province	1994	CP94017	09-AUG-1994	30.398	-81.645	1	1.0	m	
EMAP Carolinian Province	1994	CP94018	11-AUG-1994	30.516	-81.444	1	7.0	m	
EMAP Carolinian Province	1994	CP94019	11-AUG-1994	30.711	-81.47	1	8.4	m	
EMAP Carolinian Province	1994	CP94020	03-AUG-1994	30.982	-81.428	1	8.6	m	
EMAP Carolinian Province	1994	CP94021	02-AUG-1994	31.107	-81.451	1	8.5	m	
EMAP Carolinian Province	1994	CP94022	17-AUG-1994	31.391	-81.293	1	4.4	m	
EMAP Carolinian Province	1994	CP94023	15-AUG-1994	31.547	-81.19	1	5.5	m	
EMAP Carolinian Province	1994	CP94024	18-AUG-1994	31.722	-81.164	1	4.2	m	
EMAP Carolinian Province	1994	CP94025	18-AUG-1994	31.862	-81.039	1	5.5	m	
EMAP Carolinian Province	1994	CP94026	19-AUG-1994	31.93	-80.968	1	7.6	m	
EMAP Carolinian Province	1994	CP94027	25-AUG-1994	32.07	-80.919	1	4.5	m	
EMAP Carolinian Province	1994	CP94028	27-JUL-1994	33.93	-78.218	1	0.5	m	
EMAP Carolinian Province	1994	CP94029	26-JUL-1994	34.38	-77.618	1	0.5	m	
EMAP Carolinian Province	1994	CP94030	19-JUL-1994	34.506	-77.407	1	0.5	m	
EMAP Carolinian Province	1994	CP94031	01-JUL-1994	34.669	-77.152	1	0.9	m	
EMAP Carolinian Province	1994	CP94032	28-JUL-1994	34.684	-76.557	1	1.3	m	
EMAP Carolinian Province	1994	CP94033	28-JUL-1994	34.773	-76.453	1	2.0	m	
EMAP Carolinian Province	1994	CP94034	06-JUL-1994	34.973	-76.696	1	4.0	m	
EMAP Carolinian Province	1994	CP94035	06-JUL-1994	35.006	-76.408	1	3.3	m	
EMAP Carolinian Province	1994	CP94036	23-AUG-1994	35.073	-76.551	1	5.6	m	
EMAP Carolinian Province	1994	CP94037	10-AUG-1994	35.083	-76.19	1	4.6	m	
EMAP Carolinian Province	1994	CP94038	07-JUL-1994	35.096	-76.6	1	2.0	m	
EMAP Carolinian Province	1994	CP94039	10-AUG-1994	35.12	-76.028	1	2.4	m	
EMAP Carolinian Province	1994	CP94040	23-AUG-1994	35.14	-76.47	1	6.1	m	
EMAP Carolinian Province	1994	CP94041	10-AUG-1994	35.151	-76.22	1	5.9	m	
EMAP Carolinian Province	1994	CP94042	10-AUG-1994	35.16	-75.984	1	3.8	m	
EMAP Carolinian Province	1994	CP94043	23-AUG-1994	35.231	-76.56	1	2.5	m	
EMAP Carolinian Province	1994	CP94044	09-AUG-1994	35.257	-75.752	1	2.5	m	
EMAP Carolinian Province	1994	CP94045	09-AUG-1994	35.306	-75.567	1	2.3	m	
EMAP Carolinian Province	1994	CP94046	17-AUG-1994	35.343	-76.176	1	2.5	m	
EMAP Carolinian Province	1994	CP94047	16-AUG-1994	35.355	-76.694	1	3.2	m	
EMAP Carolinian Province	1994	CP94048	18-AUG-1994	35.357	-76.477	1	5.7	m	
EMAP Carolinian Province	1994	CP94049	17-AUG-1994	35.367	-76.342	1	1.7	m	
EMAP Carolinian Province	1994	CP94050	18-AUG-1994	35.379	-75.876	1	5.4	m	
EMAP Carolinian Province	1994	CP94051	16-AUG-1994	35.396	-76.675	1	4.6	m	
EMAP Carolinian Province	1994	CP94052	16-AUG-1994	35.398	-76.692	1	4.8	m	
EMAP Carolinian Province	1994	CP94053	16-AUG-1994	35.458	-76.817	1	2.7	m	
EMAP Carolinian Province	1994	CP94054	19-AUG-1994	35.476	-76.539	1	1.9	m	
EMAP Carolinian Province	1994	CP94055	02-AUG-1994	35.541	-75.716	1	4.1	m	
EMAP Carolinian Province	1994	CP94056	08-AUG-1994	35.558	-75.579	1	4.3	m	
EMAP Carolinian Province	1994	CP94057	02-AUG-1994	35.58	-75.85	1	1.3	m	
EMAP Carolinian Province	1994	CP94058	07-AUG-1994	35.657	-75.602	1	3.9	m	
EMAP Carolinian Province	1994	CP94059	08-AUG-1994	35.718	-75.564	1	1.0	m	
EMAP Carolinian Province	1994	CP94060	06-AUG-1994	35.857	-75.668	1	3.2	m	
EMAP Carolinian Province	1994	CP94061	17-JUL-1994	35.961	-76.352	1	4.0	m	
EMAP Carolinian Province	1994	CP94062	16-JUL-1994	35.991	-76.523	1	6.0	m	
EMAP Carolinian Province	1994	CP94063	16-JUL-1994	36.006	-76.536	1	1.2	m	
EMAP Carolinian Province	1994	CP94064	15-JUL-1994	36.02	-75.926	1	5.7	m	
EMAP Carolinian Province	1994	CP94065	15-JUL-1994	36.045	-76.619	1	2.5	m	
EMAP Carolinian Province	1994	CP94066	17-JUL-1994	36.053	-76.309	1	6.1	m	
EMAP Carolinian Province	1994	CP94067	17-JUL-1994	36.084	-76.456	1	2.0	m	
EMAP Carolinian Province	1994	CP94068	14-JUL-1994	36.098	-75.78	1	1.7	m	
EMAP Carolinian Province	1994	CP94069	15-JUL-1994	36.122	-75.939	1	5.5	m	
EMAP Carolinian Province	1994	CP94070	14-JUL-1994	36.145	-75.748	1	0.5	m	
EMAP Carolinian Province	1994	CP94071	13-JUL-1994	36.386	-75.855	1	0.8	m	
EMAP Carolinian Province	1994	CP94072	12-JUL-1994	36.514	-76.041	1	1.5	m	
EMAP Carolinian Province	1994	CP94073	25-AUG-1994	32.17	-80.796	1	12.9	m	
EMAP Carolinian Province	1994	CP94074	24-AUG-1994	32.28	-80.593	1	4.1	m	
EMAP Carolinian Province	1994	CP94075	23-AUG-1994	32.285	-80.749	1	10.9	m	
EMAP Carolinian Province	1994	CP94076	11-AUG-1994	32.539	-80.35	1	7.9	m	
EMAP Carolinian Province	1994	CP94077	12-AUG-1994	32.559	-80.547	1	7.5	m	
EMAP Carolinian Province	1994	CP94078	08-AUG-1994	32.614	-80.166	1	6.1	m	
EMAP Carolinian Province	1994	CP94079	29-JUL-1994	32.765	-79.887	1	10.9	m	
EMAP Carolinian Province	1994	CP94080	29-JUL-1994	32.828	-79.739	1	3.7	m	
EMAP Carolinian Province	1994	CP94081	26-JUL-1994	32.993	-79.559	1	1.2	m	
EMAP Carolinian Province	1994	CP94082	10-AUG-1994	33.359	-79.292	1	4.7	m	
EMAP Carolinian Province	1994	CP94083	29-AUG-1994	33.855	-78.565	1	5.5	m	
EMAP Carolinian Province	1994	CP94084	12-JUL-1994	36.724	-76.188	1	0.7	m	
EMAP Carolinian Province	1994	CP94CF_	29-AUG-1994	34.124	-77.927	1	2.5	m	
EMAP Carolinian Province	1994	CP94DSL	20-SEP-1994	32.816	-79.963	1	1.2	m	
EMAP Carolinian Province	1994	CP94ES4	13-JUL-1994	36.393	-75.849	1	1.0	m	
EMAP Carolinian Province	1994	CP94JAC	09-AUG-1994	30.383	-81.45	1	12.9	m	
EMAP Carolinian Province	1994	CP94KOP	03-AUG-1994	32.819	-79.964	1			
EMAP Carolinian Province	1994	CP94LTH	23-SEP-1994	32.703	-79.92	1	2.0	m	
EMAP Carolinian Province	1994	CP94MI_	26-JUL-1994	34.155	-77.85	1	2.2	m	
EMAP Carolinian Province	1994	CP94NMK	20-SEP-1994	32.807	-79.935	1	1.7	m	
EMAP Carolinian Province	1994	CP94NOI	03-AUG-1994	32.872	-79.971	1			
EMAP Carolinian Province	1994	CP94PLM	22-SEP-1994	32.763	-79.948	1	1.8	m	
EMAP Carolinian Province	1994	CP94RC_	28-JUL-1994	34.703	-76.621	1	1.6	m	
EMAP Carolinian Province	1994	CP94SPY	03-AUG-1994	32.84	-79.945	1			
EMAP Carolinian Province	1994	CP94ZI_	25-JUL-1994	33.953	-77.938	1	1.2	m	
EMAP Carolinian Province	1995	CP95101	09-AUG-1995	36.621	-75.959	1	1.4	m	
EMAP Carolinian Province	1995	CP95102	09-AUG-1995	36.421	-75.986	1	1.1	m	
EMAP Carolinian Province	1995	CP95103	08-AUG-1995	36.274	-76.689	1	3.6	m	
EMAP Carolinian Province	1995	CP95104	10-AUG-1995	36.167	-76.249	1	2.0	m	
EMAP Carolinian Province	1995	CP95105	11-AUG-1995	36.076	-75.773	1	2.2	m	
EMAP Carolinian Province	1995	CP95106	11-AUG-1995	36.041	-75.715	1	1.7	m	
EMAP Carolinian Province	1995	CP95107	10-AUG-1995	36.039	-76.269	1	6.3	m	
EMAP Carolinian Province	1995	CP95108	08-AUG-1995	35.94	-76.618	1	1.0	m	
EMAP Carolinian Province	1995	CP95109	12-AUG-1995	35.937	-76.102	1	2.2	m	
EMAP Carolinian Province	1995	CP95110	12-AUG-1995	35.917	-76.076	1	1.3	m	
EMAP Carolinian Province	1995	CP95111	12-AUG-1995	35.893	-75.88	1	1.5	m	
EMAP Carolinian Province	1995	CP95112	13-AUG-1995	35.831	-75.67	1	1.0	m	
EMAP Carolinian Province	1995	CP95113	13-AUG-1995	35.731	-75.68	1	3.8	m	
EMAP Carolinian Province	1995	CP95114	21-JUL-1995	35.514	-76.64	1	2.0	m	
EMAP Carolinian Province	1995	CP95115	25-JUL-1995	35.465	-75.575	1	4.4	m	
EMAP Carolinian Province	1995	CP95116	19-JUL-1995	35.449	-76.589	1	3.6	m	
EMAP Carolinian Province	1995	CP95117	22-JUL-1995	35.431	-75.791	1	6.0	m	
EMAP Carolinian Province	1995	CP95118	12-JUL-1995	35.422	-76.04	1	1.5	m	
EMAP Carolinian Province	1995	CP95119	12-JUL-1995	35.404	-75.943	1	5.0	m	
EMAP Carolinian Province	1995	CP95120	20-JUL-1995	35.379	-76.825	1	1.5	m	
EMAP Carolinian Province	1995	CP95121	20-JUL-1995	35.375	-76.689	1	3.8	m	
EMAP Carolinian Province	1995	CP95122	20-JUL-1995	35.372	-76.671	1	4.0	m	
EMAP Carolinian Province	1995	CP95123	26-JUL-1995	35.367	-75.611	1	4.5	m	
EMAP Carolinian Province	1995	CP95124	19-JUL-1995	35.358	-76.545	1	5.0	m	
EMAP Carolinian Province	1995	CP95125	11-JUL-1995	35.351	-76.089	1	2.5	m	
EMAP Carolinian Province	1995	CP95126	11-JUL-1995	35.34	-76.252	1	1.6	m	
EMAP Carolinian Province	1995	CP95127	11-JUL-1995	35.334	-76.305	1	2.4	m	
EMAP Carolinian Province	1995	CP95128	19-JUL-1995	35.299	-76.49	1	2.0	m	
EMAP Carolinian Province	1995	CP95129	19-JUL-1995	35.279	-76.491	1	1.0	m	
EMAP Carolinian Province	1995	CP95130	27-JUL-1995	35.273	-75.887	1	5.3	m	
EMAP Carolinian Province	1995	CP95131	29-JUL-1995	35.225	-76.152	1	6.3	m	
EMAP Carolinian Province	1995	CP95132	24-JUL-1995	35.22	-75.853	1	4.0	m	
EMAP Carolinian Province	1995	CP95133	24-JUL-1995	35.193	-75.779	1	2.3	m	
EMAP Carolinian Province	1995	CP95134	21-JUL-1995	35.148	-76.59	1	1.0	m	
EMAP Carolinian Province	1995	CP95135	23-JUL-1995	35.082	-76.003	1	0.9	m	
EMAP Carolinian Province	1995	CP95136	14-AUG-1995	35.055	-76.505	1	6.4	m	
EMAP Carolinian Province	1995	CP95138	23-AUG-1995	35.154	-76.6	1	0.8	m	
EMAP Carolinian Province	1995	CP95139	21-AUG-1995	35.009	-76.675	1	6.6	m	
EMAP Carolinian Province	1995	CP95140	21-AUG-1995	34.922	-76.661	1	1.9	m	
EMAP Carolinian Province	1995	CP95141	02-AUG-1995	34.916	-76.336	1	1.7	m	
EMAP Carolinian Province	1995	CP95142	01-AUG-1995	34.77	-76.685	1	1.3	m	
EMAP Carolinian Province	1995	CP95143	02-AUG-1995	34.754	-76.496	1	1.5	m	
EMAP Carolinian Province	1995	CP95144	31-JUL-1995	34.692	-77.106	1	0.5	m	
EMAP Carolinian Province	1995	CP95145	31-JUL-1995	34.479	-77.473	1	0.5	m	
EMAP Carolinian Province	1995	CP95146	06-JUL-1995	33.938	-77.981	1	13.0	m	
EMAP Carolinian Province	1995	CP95147	06-JUL-1995	34.034	-77.939	1	6.1	m	
EMAP Carolinian Province	1995	CP95148	05-JUL-1995	33.919	-78.372	1	2.7	m	
EMAP Carolinian Province	1995	CP95149	18-AUG-1995	33.341	-79.274	1	6.0	m	
EMAP Carolinian Province	1995	CP95150	18-AUG-1995	33.155	-79.354	1	4.2	m	
EMAP Carolinian Province	1995	CP95151	02-AUG-1995	32.785	-79.966	1	7.4	m	
EMAP Carolinian Province	1995	CP95152	02-AUG-1995	32.784	-79.962	1	9.0	m	
EMAP Carolinian Province	1995	CP95153	03-AUG-1995	32.783	-79.804	1	3.2	m	
EMAP Carolinian Province	1995	CP95154	04-AUG-1995	32.732	-79.882	1	1.2	m	
EMAP Carolinian Province	1995	CP95155	31-JUL-1995	32.602	-80.237	1	11.4	m	
EMAP Carolinian Province	1995	CP95156	01-AUG-1995	32.591	-80.398	1	6.7	m	
EMAP Carolinian Province	1995	CP95157	16-AUG-1995	32.533	-80.572	1	10.6	m	
EMAP Carolinian Province	1995	CP95158	15-AUG-1995	32.512	-80.606	1	4.8	m	
EMAP Carolinian Province	1995	CP95159	28-AUG-1995	32.266	-80.694	1	11.1	m	
EMAP Carolinian Province	1995	CP95160	29-AUG-1995	32.248	-80.753	1	2.1	m	
EMAP Carolinian Province	1995	CP95161	30-AUG-1995	32.08	-80.88	1	5.3	m	
EMAP Carolinian Province	1995	CP95162	29-AUG-1995	32.026	-80.912	1	3.6	m	
EMAP Carolinian Province	1995	CP95163	29-AUG-1995	31.986	-80.929	1	8.4	m	
EMAP Carolinian Province	1995	CP95164	22-AUG-1995	31.861	-81.109	1	6.6	m	
EMAP Carolinian Province	1995	CP95165	08-SEP-1995	31.689	-81.192	1	8.0	m	
EMAP Carolinian Province	1995	CP95166	07-SEP-1995	31.494	-81.294	1	2.1	m	
EMAP Carolinian Province	1995	CP95167	05-SEP-1995	31.257	-81.326	1	3.5	m	
EMAP Carolinian Province	1995	CP95168	06-SEP-1995	31.072	-81.495	1	7.1	m	
EMAP Carolinian Province	1995	CP95169	07-SEP-1995	30.927	-81.462	1	6.1	m	
EMAP Carolinian Province	1995	CP95170	04-AUG-1995	30.559	-81.47	1	5.0	m	
EMAP Carolinian Province	1995	CP95171	03-AUG-1995	30.393	-81.554	1	11.0	m	
EMAP Carolinian Province	1995	CP95172	16-AUG-1995	30.135	-81.731	1	3.0	m	
EMAP Carolinian Province	1995	CP95173	08-AUG-1995	29.564	-81.185	1	5.0	m	
EMAP Carolinian Province	1995	CP95174	07-AUG-1995	29.24	-81.027	1	1.5	m	
EMAP Carolinian Province	1995	CP95175	09-AUG-1995	28.74	-80.796	1	1.6	m	
EMAP Carolinian Province	1995	CP95176	31-JUL-1995	28.502	-80.749	1	1.5	m	
EMAP Carolinian Province	1995	CP95177	31-JUL-1995	28.464	-80.739	1	1.7	m	
EMAP Carolinian Province	1995	CP95178	27-JUL-1995	28.368	-80.681	1	1.3	m	
EMAP Carolinian Province	1995	CP95179	26-JUL-1995	28.353	-80.674	1	0.9	m	
EMAP Carolinian Province	1995	CP95180	25-JUL-1995	28.293	-80.685	1	2.2	m	
EMAP Carolinian Province	1995	CP95181	24-JUL-1995	28.142	-80.618	1	3.4	m	
EMAP Carolinian Province	1995	CP95182	10-AUG-1995	27.994	-80.535	1	2.0	m	
EMAP Carolinian Province	1995	CP95183	18-AUG-1995	27.827	-80.451	1	1.6	m	
EMAP Carolinian Province	1995	CP95184	21-AUG-1995	27.714	-80.4	1	0.6	m	
EMAP Carolinian Province	1995	CP95185	22-AUG-1995	27.578	-80.357	1	1.3	m	
EMAP Carolinian Province	1995	CP95186	23-AUG-1995	27.365	-80.266	1	1.6	m	
EMAP Carolinian Province	1995	CP95187	23-AUG-1995	27.346	-80.268	1	2.0	m	
EMAP Carolinian Province	1995	CP95188	25-AUG-1995	27.271	-80.222	1	2.3	m	
EMAP Carolinian Province	1995	CP95ASM	27-SEP-1995	32.78	-79.955	1	0.8	m	
EMAP Carolinian Province	1995	CP95CB_	11-AUG-1995	36.4	-75.845	1	1.0	m	
EMAP Carolinian Province	1995	CP95CF_	22-AUG-1995	34.124	-77.927	1	1.4	m	
EMAP Carolinian Province	1995	CP95DIE	26-SEP-1995	32.804	-79.966	1	1.2	m	
EMAP Carolinian Province	1995	CP95FOS	10-OCT-1995	32.86	-79.855	1	2.5	m	
EMAP Carolinian Province	1995	CP95KIA	12-OCT-1995	32.603	-80.132	1			
EMAP Carolinian Province	1995	CP95KOP	26-SEP-1995	32.829	-79.965	1	1.7	m	
EMAP Carolinian Province	1995	CP95LON	12-OCT-1995	32.685	-80.123	1			
EMAP Carolinian Province	1995	CP95LTH	25-OCT-1995	32.702	-79.92	1	2.4	m	
EMAP Carolinian Province	1995	CP95MI_	03-AUG-1995	34.156	-77.85	1	0.9	m	
EMAP Carolinian Province	1995	CP95NMK	06-OCT-1995	32.807	-79.941	1	1.7	m	
EMAP Carolinian Province	1995	CP95NV1	04-OCT-1995	32.867	-79.964	1	8.1	m	
EMAP Carolinian Province	1995	CP95NV2	04-OCT-1995	32.846	-79.933	1	3.0	m	
EMAP Carolinian Province	1995	CP95PR1	14-SEP-1995	35.354	-76.653	1	2.9	m	
EMAP Carolinian Province	1995	CP95PR2	14-SEP-1995	35.368	-76.617	1	4.8	m	
EMAP Carolinian Province	1995	CP95PR3	14-SEP-1995	35.401	-76.751	1	4.6	m	
EMAP Carolinian Province	1995	CP95PR4	14-SEP-1995	35.408	-76.775	1	4.0	m	
EMAP Carolinian Province	1995	CP95PR5	14-SEP-1995	35.434	-76.826	1	4.3	m	
EMAP Carolinian Province	1995	CP95RC_	01-AUG-1995	34.711	-76.647	1	0.5	m	
EMAP Carolinian Province	1995	CP95SPY	27-SEP-1995	32.839	-79.945	1	2.5	m	
EMAP Carolinian Province	1995	CP95ZI_	22-AUG-1995	33.956	-77.939	1	1.0	m	
EMAP Carolinian Province	1996	CP96201	19-SEP-1996	36.495	-76.005	1	2.1	m	
EMAP Carolinian Province	1996	CP96202	18-SEP-1996	36.281	-76.151	1	3.6	m	
EMAP Carolinian Province	1996	CP96203	18-SEP-1996	36.237	-75.81	1	1.0	m	
EMAP Carolinian Province	1996	CP96204	18-SEP-1996	36.155	-75.796	1	3.0	m	
EMAP Carolinian Province	1996	CP96205	09-JUL-1996	36.13	-76.333	1	3.5	m	
EMAP Carolinian Province	1996	CP96206	17-SEP-1996	36.104	-75.954	1	5.6	m	
EMAP Carolinian Province	1996	CP96207	09-JUL-1996	36.069	-76.274	1	6.2	m	
EMAP Carolinian Province	1996	CP96208	19-SEP-1996	35.952	-75.661	1	2.7	m	
EMAP Carolinian Province	1996	CP96209	19-SEP-1996	35.944	-75.885	1	2.3	m	
EMAP Carolinian Province	1996	CP96210	10-JUL-1996	35.936	-76.302	1	3.1	m	
EMAP Carolinian Province	1996	CP96211	10-JUL-1996	35.93	-76.736	1	2.7	m	
EMAP Carolinian Province	1996	CP96212	19-SEP-1996	35.828	-75.684	1	3.5	m	
EMAP Carolinian Province	1996	CP96213	19-SEP-1996	35.733	-75.642	1	4.4	m	
EMAP Carolinian Province	1996	CP96214	10-JUL-1996	35.542	-76.632	1	1.4	m	
EMAP Carolinian Province	1996	CP96215	16-SEP-1996	35.511	-75.967	1	1.8	m	
EMAP Carolinian Province	1996	CP96216	16-SEP-1996	35.46	-75.579	1	4.8	m	
EMAP Carolinian Province	1996	CP96217	22-JUL-1996	35.43	-76.667	1	0.9	m	
EMAP Carolinian Province	1996	CP96218	16-SEP-1996	35.417	-75.788	1	6.4	m	
EMAP Carolinian Province	1996	CP96219	16-SEP-1996	35.404	-75.945	1	5.2	m	
EMAP Carolinian Province	1996	CP96220	23-JUL-1996	35.395	-76.416	1	2.6	m	
EMAP Carolinian Province	1996	CP96221	22-JUL-1996	35.389	-76.669	1	4.2	m	
EMAP Carolinian Province	1996	CP96222	16-SEP-1996	35.372	-75.609	1	5.0	m	
EMAP Carolinian Province	1996	CP96223	23-JUL-1996	35.34	-76.287	1	1.6	m	
EMAP Carolinian Province	1996	CP96224	16-SEP-1996	35.339	-76.088	1	2.3	m	
EMAP Carolinian Province	1996	CP96225	22-JUL-1996	35.335	-76.5	1	4.5	m	
EMAP Carolinian Province	1996	CP96226	22-JUL-1996	35.332	-76.612	1	1.5	m	
EMAP Carolinian Province	1996	CP96227	16-SEP-1996	35.275	-75.889	1	6.1	m	
EMAP Carolinian Province	1996	CP96228	23-JUL-1996	35.263	-76.476	1	0.9	m	
EMAP Carolinian Province	1996	CP96229	16-SEP-1996	35.235	-75.85	1	4.6	m	
EMAP Carolinian Province	1996	CP96230	15-SEP-1996	35.235	-76.152	1	6.2	m	
EMAP Carolinian Province	1996	CP96231	16-SEP-1996	35.192	-75.78	1	0.6	m	
EMAP Carolinian Province	1996	CP96232	25-JUL-1996	35.168	-76.667	1	3.5	m	
EMAP Carolinian Province	1996	CP96233	24-JUL-1996	35.085	-76.519	1	6.8	m	
EMAP Carolinian Province	1996	CP96234	16-SEP-1996	35.081	-76.024	1	1.4	m	
EMAP Carolinian Province	1996	CP96235	24-JUL-1996	35.002	-76.689	1	5.7	m	
EMAP Carolinian Province	1996	CP96236	24-JUL-1996	34.991	-76.5	1	1.4	m	
EMAP Carolinian Province	1996	CP96237	12-SEP-1996	34.862	-76.403	1	2.6	m	
EMAP Carolinian Province	1996	CP96238	25-JUL-1996	34.705	-76.912	1	1.0	m	
EMAP Carolinian Province	1996	CP96239	13-SEP-1996	34.625	-76.537	1	3.6	m	
EMAP Carolinian Province	1996	CP96240	25-JUL-1996	34.566	-77.365	1	1.2	m	
EMAP Carolinian Province	1996	CP96241	29-JUL-1996	34.133	-77.865	1	1.2	m	
EMAP Carolinian Province	1996	CP96242	29-JUL-1996	34.109	-77.867	1	0.1	m	
EMAP Carolinian Province	1997	CP97022	14-AUG-1997	31.391	-81.293	1	3.8	m	
EMAP Carolinian Province	1997	CP97036	17-JUL-1997	35.073	-76.551	1	5.2	m	
EMAP Carolinian Province	1997	CP97052	15-JUL-1997	35.398	-76.692	1	4.4	m	
EMAP Carolinian Province	1997	CP97071	23-AUG-1997	36.386	-75.855	1	1.0	m	
EMAP Carolinian Province	1997	CP97075	30-JUL-1997	32.285	-80.749	1	9.9	m	
EMAP Carolinian Province	1997	CP97082	24-JUL-1997	33.359	-79.292	1	4.6	m	
EMAP Carolinian Province	1997	CP97109	08-JUL-1997	35.937	-76.102	1	2.6	m	
EMAP Carolinian Province	1997	CP97114	16-JUL-1997	35.514	-76.64	1	2.0	m	
EMAP Carolinian Province	1997	CP97120	15-JUL-1997	35.379	-76.825	1	1.4	m	
EMAP Carolinian Province	1997	CP97141	23-JUL-1997	34.916	-76.336	1	2.0	m	
EMAP Carolinian Province	1997	CP97149	24-JUL-1997	33.341	-79.274	1	4.7	m	
EMAP Carolinian Province	1997	CP97156	22-JUL-1997	32.591	-80.398	1	8.2	m	
EMAP Carolinian Province	1997	CP97164	29-JUL-1997	31.861	-81.109	1	6.7	m	
EMAP Carolinian Province	1997	CP97172	13-AUG-1997	30.135	-81.731	1	3.1	m	
EMAP Carolinian Province	1997	CP97183	12-AUG-1997	27.827	-80.451	1			
EMAP Carolinian Province	1997	CP97184	12-AUG-1997	27.714	-80.4	1			
EMAP Carolinian Province	1997	CP97301	23-AUG-1997	36.518	-75.98	1	1.2	m	
EMAP Carolinian Province	1997	CP97302	23-AUG-1997	36.413	-75.9	1	1.0	m	
EMAP Carolinian Province	1997	CP97303	22-AUG-1997	36.235	-75.934	1	3.7	m	
EMAP Carolinian Province	1997	CP97304	23-AUG-1997	36.23	-75.816	1	1.2	m	
EMAP Carolinian Province	1997	CP97305	22-AUG-1997	36.149	-75.781	1	2.3	m	
EMAP Carolinian Province	1997	CP97306	20-AUG-1997	36.137	-76.131	1	1.0	m	
EMAP Carolinian Province	1997	CP97307	22-AUG-1997	36.087	-75.964	1	5.3	m	
EMAP Carolinian Province	1997	CP97308	20-AUG-1997	36.072	-76.275	1	5.1	m	
EMAP Carolinian Province	1997	CP97309	22-AUG-1997	35.952	-76.714	1	1.7	m	
EMAP Carolinian Province	1997	CP97310	08-JUL-1997	35.92	-75.982	1	3.6	m	
EMAP Carolinian Province	1997	CP97311	21-AUG-1997	35.917	-76.721	1	4.6	m	
EMAP Carolinian Province	1997	CP97312	08-SEP-1997	35.824	-75.677	1	4.4	m	
EMAP Carolinian Province	1997	CP97313	09-JUL-1997	35.739	-75.636	1	3.4	m	
EMAP Carolinian Province	1997	CP97314	08-JUL-1997	35.698	-75.757	1	1.2	m	
EMAP Carolinian Province	1997	CP97315	16-JUL-1997	35.5	-77.03	1	1.4	m	
EMAP Carolinian Province	1997	CP97316	19-AUG-1997	35.448	-75.587	1	5.1	m	
EMAP Carolinian Province	1997	CP97317	11-JUL-1997	35.429	-76.532	1	2.1	m	
EMAP Carolinian Province	1997	CP97318	19-AUG-1997	35.412	-75.779	1	6.0	m	
EMAP Carolinian Province	1997	CP97319	10-JUL-1997	35.406	-75.967	1	4.4	m	
EMAP Carolinian Province	1997	CP97320	15-JUL-1997	35.406	-76.752	1	4.6	m	
EMAP Carolinian Province	1997	CP97321	11-JUL-1997	35.388	-76.46	1	2.7	m	
EMAP Carolinian Province	1997	CP97322	11-JUL-1997	35.376	-76.65	1	4.6	m	
EMAP Carolinian Province	1997	CP97323	10-JUL-1997	35.359	-76.131	1	0.7	m	
EMAP Carolinian Province	1997	CP97324	19-AUG-1997	35.37	-75.583	1	4.0	m	
EMAP Carolinian Province	1997	CP97325	10-JUL-1997	35.339	-76.288	1	2.0	m	
EMAP Carolinian Province	1997	CP97326	18-AUG-1997	35.322	-76.055	1	3.4	m	
EMAP Carolinian Province	1997	CP97327	11-JUL-1997	35.321	-76.558	1	1.5	m	
EMAP Carolinian Province	1997	CP97328	19-AUG-1997	35.275	-75.88	1	5.3	m	
EMAP Carolinian Province	1997	CP97329	23-JUL-1997	35.237	-76.514	1	0.8	m	
EMAP Carolinian Province	1997	CP97330	19-AUG-1997	35.236	-76.148	1	5.4	m	
EMAP Carolinian Province	1997	CP97331	18-AUG-1997	35.233	-75.849	1	4.3	m	
EMAP Carolinian Province	1997	CP97332	19-AUG-1997	35.192	-75.765	1	3.6	m	
EMAP Carolinian Province	1997	CP97333	18-JUL-1997	35.071	-77.076	1	2.0	m	
EMAP Carolinian Province	1997	CP97334	17-JUL-1997	35.089	-76.514	1	6.6	m	
EMAP Carolinian Province	1997	CP97335	18-AUG-1997	35.077	-76.014	1	0.9	m	
EMAP Carolinian Province	1997	CP97336	17-JUL-1997	35.0	-76.684	1	5.6	m	
EMAP Carolinian Province	1997	CP97337	23-JUL-1997	34.975	-76.278	1	2.5	m	
EMAP Carolinian Province	1997	CP97338	17-JUL-1997	34.967	-76.583	1	2.9	m	
EMAP Carolinian Province	1997	CP97339	24-JUL-1997	34.761	-76.604	1	1.2	m	
EMAP Carolinian Province	1997	CP97340	22-JUL-1997	34.717	-76.562	1	3.2	m	
EMAP Carolinian Province	1997	CP97341	22-JUL-1997	34.7	-76.671	1	6.0	m	
EMAP Carolinian Province	1997	CP97342	03-JUL-1997	34.266	-77.77	1	1.3	m	
EMAP Carolinian Province	1997	CP97343	03-JUL-1997	33.9	-78.028	1	2.3	m	
EMAP Carolinian Province	1997	CP97345	21-AUG-1997	36.461	-76.996	1	9.3	m	
EMAP Carolinian Province	1997	CP97346	21-AUG-1997	36.396	-76.92	1	6.8	m	
EMAP Carolinian Province	1997	CP97347	21-AUG-1997	36.375	-76.846	1	6.4	m	
EMAP Carolinian Province	1997	CP97348	21-AUG-1997	36.363	-76.79	1	2.0	m	
EMAP Carolinian Province	1997	CP97349	21-AUG-1997	36.292	-76.698	1	3.7	m	
EMAP Carolinian Province	1997	CP97350	21-AUG-1997	36.218	-76.718	1	7.0	m	
EMAP Carolinian Province	1997	CP97351	21-AUG-1997	36.174	-76.745	1	4.5	m	
EMAP Carolinian Province	1997	CP97352	21-AUG-1997	36.117	-76.737	1	6.1	m	
EMAP Carolinian Province	1997	CP97353	21-AUG-1997	36.083	-76.718	1	5.4	m	
EMAP Carolinian Province	1997	CP97354	21-AUG-1997	36.026	-76.666	1	4.0	m	
EMAP Carolinian Province	1997	CP97HOB	31-AUG-1997	32.826	-79.873	1			
EMAP Carolinian Province	1997	CP97JIY	29-AUG-1997	32.756	-79.918	1			
EMAP Carolinian Province	1997	CP97SPY	29-AUG-1997	32.838	-79.946	1			
EMAP Carolinian Province	1997	CP97WAN	29-AUG-1997	32.811	-79.909	1			
National Coastal Assessment-Southeast/Florida Fish and Wildlife Research Institute	2000	FL00-0005	06-JUL-2000	30.425	-81.539	1	0.6	m	
National Coastal Assessment-Southeast/Florida Fish and Wildlife Research Institute	2000	FL00-0006	12-JUL-2000	30.247	-81.652	1	4.5	m	
National Coastal Assessment-Southeast/Florida Fish and Wildlife Research Institute	2000	FL00-0008	12-JUL-2000	30.209	-81.677	1	2.0	m	
National Coastal Assessment-Southeast/Florida Fish and Wildlife Research Institute	2000	FL00-0012	22-AUG-2000	28.739	-80.72	1	1.6	m	
National Coastal Assessment-Southeast/Florida Fish and Wildlife Research Institute	2000	FL00-0013	22-AUG-2000	28.426	-80.639	1	2.1	m	
National Coastal Assessment-Southeast/Florida Fish and Wildlife Research Institute	2000	FL00-0015	23-AUG-2000	27.857	-80.462	1	1.5	m	
National Coastal Assessment-Southeast/Florida Fish and Wildlife Research Institute	2001	FL01-0004	13-AUG-2001	30.376	-81.622	1	5.7	m	
National Coastal Assessment-Southeast/Florida Fish and Wildlife Research Institute	2001	FL01-0005	14-AUG-2001	30.264	-81.697	1	0.4	m	
National Coastal Assessment-Southeast/Florida Fish and Wildlife Research Institute	2001	FL01-0006	14-AUG-2001	30.102	-81.668	1	3.6	m	
National Coastal Assessment-Southeast/Florida Fish and Wildlife Research Institute	2001	FL01-0009	13-AUG-2001	30.425	-81.539	1	1.0	m	
National Coastal Assessment-Southeast/Florida Fish and Wildlife Research Institute	2001	FL01-0011	23-JUL-2001	28.427	-80.639	1	2.2	m	
National Coastal Assessment-Southeast/Florida Fish and Wildlife Research Institute	2002	FL02-0020	08-JUL-2002	28.426	-80.639	1	2.2	m	
National Coastal Assessment-Southeast/Florida Fish and Wildlife Research Institute	2002	FL02-0022	17-JUL-2002	30.425	-81.539	1	1.0	m	
National Coastal Assessment-Southeast/Florida Fish and Wildlife Research Institute	2003	FL03-0004	14-JUL-2003	28.426	-80.639	4	1.9	m	
National Coastal Assessment-Southeast/Florida Fish and Wildlife Research Institute	2003	FL03-0005	15-JUL-2003	30.425	-81.539	4	1.1	m	
National Coastal Assessment-Southeast/Florida Fish and Wildlife Research Institute	2003	FL03-0009	04-AUG-2003	28.492	-80.761	1	2.2	m	
National Coastal Assessment-Southeast/Florida Fish and Wildlife Research Institute	2004	FL04-0006	08-JUL-2004	30.567	-81.507	1			
National Coastal Assessment-Southeast/Florida Fish and Wildlife Research Institute	2004	FL04-0032	14-JUL-2004	29.34	-81.079	1	1.0	m	
National Coastal Assessment-Southeast/Florida Fish and Wildlife Research Institute	2004	FL04-0043	02-AUG-2004	27.832	-80.446	1	1.9	m	
National Coastal Assessment-Southeast/Florida Fish and Wildlife Research Institute	2004	FL04-0044	27-JUL-2004	30.257	-81.663	1			
National Coastal Assessment-Southeast/Florida Fish and Wildlife Research Institute	2004	FL04-0045	03-AUG-2004	28.407	-80.744	1	1.8	m	
National Coastal Assessment-Southeast/Florida Fish and Wildlife Research Institute	2004	FL04-0050	05-AUG-2004	30.129	-81.738	1			
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0001	01-SEP-2000	31.92	-80.965	1	2.3	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0002	31-AUG-2000	31.913	-80.915	1	8.4	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0003	28-AUG-2000	31.839	-81.05	1	4.3	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0004	11-AUG-2000	31.524	-81.29	1	5.1	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0005	11-AUG-2000	31.534	-81.229	1	2.8	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0006	06-JUL-2000	31.108	-81.425	1	7.3	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0007	13-JUL-2000	31.043	-81.463	1	5.0	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0008	25-JUL-2000	30.946	-81.435	1	6.4	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0009	26-JUL-2000	30.776	-81.47	1	4.7	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0010	26-JUL-2000	30.739	-81.479	1	4.4	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0011	01-SEP-2000	31.956	-80.933	1	4.6	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0012	11-AUG-2000	31.488	-81.323	1	5.9	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0013	08-AUG-2000	31.433	-81.294	1	7.8	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0014	13-JUL-2000	31.065	-81.526	1	3.7	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0015	25-JUL-2000	30.906	-81.464	1	3.3	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0016	25-JUL-2000	30.863	-81.497	1	7.7	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0017	28-AUG-2000	31.893	-81.205	1	2.4	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0018	28-AUG-2000	31.912	-81.135	1	6.0	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0019	23-AUG-2000	31.676	-81.216	1	6.4	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0020	23-AUG-2000	31.675	-81.255	1	3.8	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0021	23-AUG-2000	31.555	-81.23	1	3.7	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0022	08-AUG-2000	31.412	-81.301	1	4.3	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0023	05-JUL-2000	31.183	-81.525	1	10.6	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0024	21-JUL-2000	30.99	-81.418	1	5.5	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0025	25-JUL-2000	30.969	-81.505	1	7.9	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0026	26-JUL-2000	30.864	-81.579	1	2.2	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0027	30-AUG-2000	32.147	-81.141	1	3.4	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0028	30-AUG-2000	32.099	-81.01	1	2.4	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0029	30-AUG-2000	32.092	-81.023	1	6.1	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0030	01-SEP-2000	32.076	-80.987	1	2.3	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0031	01-SEP-2000	32.058	-80.948	1	2.4	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0032	30-AUG-2000	32.064	-81.025	1	2.1	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0033	29-AUG-2000	32.03	-80.99	1	0.9	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0034	25-AUG-2000	31.796	-81.148	1	3.2	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0035	25-AUG-2000	31.772	-81.202	1	0.9	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0036	24-AUG-2000	31.756	-81.247	1	3.7	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0037	24-AUG-2000	31.731	-81.197	1	4.6	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0038	24-AUG-2000	31.741	-81.22	1	2.7	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0039	24-AUG-2000	31.719	-81.154	1	2.3	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0040	11-AUG-2000	31.576	-81.314	1	4.1	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0041	08-AUG-2000	31.333	-81.386	1	2.7	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0042	12-SEP-2000	31.298	-81.285	1	1.8	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0043	11-JUL-2000	31.288	-81.379	1	3.4	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0044	11-JUL-2000	31.243	-81.422	1	4.0	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0045	11-JUL-2000	31.239	-81.325	1	6.4	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0046	11-JUL-2000	31.239	-81.422	1	3.6	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0047	06-JUL-2000	31.138	-81.421	1	7.0	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0048	13-JUL-2000	31.079	-81.531	1	2.6	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0049	21-JUL-2000	31.01	-81.455	1	1.8	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2000	GA00-0050	26-JUL-2000	30.726	-81.507	1	2.8	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0001	31-JUL-2001	30.863	-81.497	1	3.3	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0002	12-JUL-2001	30.99	-81.418	1	3.9	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0003	16-AUG-2001	31.731	-81.197	1	4.6	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0004	16-AUG-2001	31.741	-81.22	1	2.2	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0005	11-JUL-2001	31.079	-81.53	1	4.8	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0006	29-AUG-2001	32.13	-81.12	1	2.1	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0007	29-AUG-2001	32.113	-81.113	1	2.7	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0008	29-AUG-2001	32.084	-81.043	1	4.1	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0009	29-AUG-2001	32.076	-80.994	1	4.2	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0010	27-AUG-2001	32.021	-80.99	1	2.7	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0011	27-AUG-2001	31.997	-81.004	1	1.5	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0012	24-AUG-2001	31.979	-81.291	1	3.3	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0013	22-AUG-2001	31.93	-81.276	1	3.4	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0014	22-AUG-2001	31.902	-81.198	1	2.2	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0015	16-AUG-2001	31.841	-81.336	1	1.8	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0016	17-AUG-2001	31.748	-81.158	1	1.6	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0017	17-AUG-2001	31.732	-81.159	1	1.2	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0018	17-AUG-2001	31.707	-81.142	1	7.0	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0019	08-AUG-2001	31.544	-81.321	1	2.5	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0020	08-AUG-2001	31.517	-81.262	1	1.7	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0021	09-AUG-2001	31.333	-81.343	1	2.7	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0022	02-AUG-2001	31.313	-81.296	1	1.4	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0023	09-AUG-2001	31.321	-81.341	1	3.2	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0024	13-JUL-2001	31.316	-81.437	1	4.0	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0025	09-AUG-2001	31.31	-81.389	1	2.0	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0026	02-AUG-2001	31.304	-81.308	1	1.8	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0027	10-JUL-2001	31.182	-81.461	1	4.8	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0028	03-JUL-2001	31.177	-81.708	1	1.4	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0029	11-JUL-2001	31.109	-81.531	1	1.2	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0030	10-JUL-2001	31.068	-81.43	1	1.2	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0031	11-JUL-2001	31.043	-81.457	1	4.8	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0032	11-JUL-2001	31.029	-81.481	1	3.4	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0033	28-AUG-2001	31.979	-80.984	1	3.4	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0034	30-AUG-2001	31.928	-80.961	1	2.6	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0035	23-AUG-2001	31.857	-81.013	1	6.1	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0036	23-AUG-2001	31.853	-81.052	1	2.4	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0037	23-AUG-2001	31.836	-81.032	1	3.7	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0038	23-AUG-2001	31.786	-81.104	1	4.5	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0039	16-AUG-2001	31.695	-81.182	1	7.4	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0040	14-AUG-2001	31.692	-81.202	1	3.4	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0041	08-AUG-2001	31.544	-81.19	1	13.5	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0042	03-JUL-2001	31.216	-81.879	1	4.1	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0043	03-JUL-2001	31.191	-81.823	1	1.8	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0044	19-JUL-2001	30.988	-81.519	1	2.9	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0045	12-JUL-2001	30.973	-81.492	1	6.1	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0046	19-JUL-2001	30.913	-81.519	1	1.8	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0047	31-JUL-2001	30.856	-81.579	1	1.8	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0048	20-JUL-2001	30.826	-81.504	1	5.9	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0049	31-JUL-2001	30.774	-81.475	1	2.0	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2001	GA01-0050	31-JUL-2001	30.759	-81.48	1	0.9	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0001	10-JUL-2002	30.862	-81.497	1	5.9	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0002	17-JUL-2002	30.99	-81.418	1	3.8	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0003	06-AUG-2002	31.73	-81.197	1	5.4	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0004	06-AUG-2002	31.74	-81.219	1	4.0	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0005	18-JUL-2002	31.078	-81.53	1	5.2	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0006	27-AUG-2002	32.085	-81.048	1	3.6	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0007	28-AUG-2002	32.037	-80.961	1	4.6	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0008	27-AUG-2002	32.04	-80.909	1	1.5	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0009	20-AUG-2002	31.991	-81.004	1	1.8	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0010	20-AUG-2002	31.977	-81.044	1	1.7	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0011	28-AUG-2002	31.983	-80.911	1	1.5	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0012	20-AUG-2002	31.979	-81.006	1	3.5	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0013	13-AUG-2002	31.908	-81.263	1	3.0	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0014	14-AUG-2002	31.864	-81.103	1	2.3	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0015	07-AUG-2002	31.825	-81.347	1	1.2	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0016	07-AUG-2002	31.819	-81.314	1	2.6	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0017	06-AUG-2002	31.794	-81.165	1	4.4	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0018	06-AUG-2002	31.737	-81.155	1	4.8	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0019	06-AUG-2002	31.726	-81.147	1	7.2	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0020	01-AUG-2002	31.528	-81.285	1	0.8	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0021	30-JUL-2002	31.49	-81.302	1	1.7	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0022	24-JUL-2002	31.312	-81.297	1	1.2	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0023	24-JUL-2002	31.309	-81.28	1	0.9	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0024	23-JUL-2002	31.273	-81.387	1	1.2	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0025	23-JUL-2002	31.182	-81.361	1	2.0	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0026	08-AUG-2002	31.134	-81.42	1	8.0	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0027	21-AUG-2002	31.122	-81.404	1	2.6	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0028	08-AUG-2002	31.113	-81.428	1	11.2	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0029	18-JUL-2002	31.056	-81.526	1	1.1	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0030	18-JUL-2002	31.033	-81.444	1	2.7	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0031	09-JUL-2002	30.733	-81.573	1	4.9	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0032	10-JUL-2002	30.725	-81.503	1	3.0	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0033	20-AUG-2002	31.941	-81.08	1	1.5	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0034	28-AUG-2002	31.916	-80.972	1	1.5	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0035	14-AUG-2002	31.928	-81.173	1	1.4	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0036	14-AUG-2002	31.852	-81.048	1	2.7	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0037	14-AUG-2002	31.851	-81.019	1	3.4	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0038	01-AUG-2002	31.574	-81.223	1	5.6	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0039	01-AUG-2002	31.556	-81.258	1	2.4	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0040	26-JUL-2002	31.473	-81.292	1	1.2	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0041	26-JUL-2002	31.449	-81.338	1	7.0	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0042	26-JUL-2002	31.347	-81.286	1	1.2	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0043	17-JUL-2002	31.0	-81.459	1	1.2	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0044	17-JUL-2002	30.978	-81.576	1	3.9	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0045	17-JUL-2002	30.965	-81.486	1	1.2	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0046	17-JUL-2002	30.96	-81.433	1	5.9	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0047	11-JUL-2002	30.905	-81.458	1	2.3	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0048	11-JUL-2002	30.884	-81.541	1	1.2	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0049	10-JUL-2002	30.844	-81.476	1	1.2	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2002	GA02-0050	09-JUL-2002	30.768	-81.488	1	8.5	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0001	10-JUL-2003	30.863	-81.497	1	7.0	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0002	09-JUL-2003	30.984	-81.42	1	11.9	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0003	06-AUG-2003	31.731	-81.197	1	6.3	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0004	06-AUG-2003	31.741	-81.219	1	3.0	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0005	15-JUL-2003	31.079	-81.53	1	7.2	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0006	27-AUG-2003	32.107	-80.999	1	5.0	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0007	27-AUG-2003	32.101	-81.085	1	0.5	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0008	28-AUG-2003	32.069	-80.976	1	3.9	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0009	27-AUG-2003	32.087	-81.064	1	0.8	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0010	28-AUG-2003	32.039	-80.981	1	2.3	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0011	28-AUG-2003	31.993	-80.938	1	3.7	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0012	21-AUG-2003	31.979	-81.046	1	5.5	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0013	13-AUG-2003	31.979	-81.292	1	3.7	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0014	19-AUG-2003	31.852	-81.104	1	0.8	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0015	14-AUG-2003	31.839	-81.154	1	7.3	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0016	14-AUG-2003	31.815	-81.143	1	3.7	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0017	12-AUG-2003	31.776	-81.277	1	5.4	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0018	07-AUG-2003	31.744	-81.161	1	7.2	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0019	07-AUG-2003	31.713	-81.166	1	3.2	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0020	07-AUG-2003	31.701	-81.146	1	7.9	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0021	30-JUL-2003	31.564	-81.356	1	2.7	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0022	30-JUL-2003	31.531	-81.353	1	1.2	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0023	29-JUL-2003	31.333	-81.355	1	2.2	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0024	22-JUL-2003	31.33	-81.32	1	0.8	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0025	29-JUL-2003	31.302	-81.288	1	0.6	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0026	31-JUL-2003	31.315	-81.377	1	0.8	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0027	22-JUL-2003	31.211	-81.437	1	2.5	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0028	29-JUL-2003	31.207	-81.342	1	0.8	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0029	08-JUL-2003	31.106	-81.451	1	7.9	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0030	15-JUL-2003	31.098	-81.551	1	3.7	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0031	15-JUL-2003	31.057	-81.501	1	6.2	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0032	09-JUL-2003	31.024	-81.446	1	2.5	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0033	21-AUG-2003	31.953	-80.929	1	1.1	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0034	20-AUG-2003	31.935	-81.158	1	7.7	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0035	20-AUG-2003	31.893	-81.103	1	1.7	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0036	19-AUG-2003	31.852	-81.041	1	1.7	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0037	12-AUG-2003	31.668	-81.265	1	6.6	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0038	30-JUL-2003	31.605	-81.247	1	3.8	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0039	24-JUL-2003	31.549	-81.181	1	5.5	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0040	23-JUL-2003	31.45	-81.355	1	1.4	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0041	23-JUL-2003	31.412	-81.352	1	1.8	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0042	23-JUL-2003	31.419	-81.306	1	0.9	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0043	22-JUL-2003	31.359	-81.372	1	1.9	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0044	08-JUL-2003	31.21	-81.596	1	3.3	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0045	07-JUL-2003	31.111	-81.481	1	7.0	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0046	09-JUL-2003	30.999	-81.457	1	1.1	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0047	18-JUL-2003	30.902	-81.457	1	6.3	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0048	10-JUL-2003	30.863	-81.563	1	3.0	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0049	10-JUL-2003	30.816	-81.496	1	3.6	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2003	GA03-0050	10-JUL-2003	30.762	-81.476	1	0.9	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0001	14-JUL-2004	30.858	-81.492	1	5.2	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0002	24-JUN-2004	30.984	-81.419	1	12.9	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0003	28-JUL-2004	31.725	-81.192	1	3.9	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0004	28-JUL-2004	31.738	-81.218	1	1.6	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0005	01-JUL-2004	31.074	-81.524	1	6.6	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0006	12-AUG-2004	32.168	-81.136	1	1.5	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0007	12-AUG-2004	32.093	-81.003	1	0.9	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0008	19-AUG-2004	32.07	-80.97	1	5.1	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0009	19-AUG-2004	32.006	-81.007	1	1.5	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0010	19-AUG-2004	31.951	-80.986	1	1.2	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0011	04-AUG-2004	31.9	-81.176	1	2.1	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0012	05-AUG-2004	31.887	-81.217	1	1.2	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0013	28-JUL-2004	31.81	-81.308	1	1.6	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0014	04-AUG-2004	31.771	-81.193	1	4.7	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0015	29-JUL-2004	31.752	-81.17	1	8.4	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0016	29-JUL-2004	31.704	-81.157	1	9.1	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0017	21-JUL-2004	31.543	-81.326	1	9.8	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0018	21-JUL-2004	31.535	-81.357	1	3.7	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0019	21-JUL-2004	31.536	-81.287	1	3.7	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0020	22-JUL-2004	31.51	-81.256	1	5.2	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0021	13-JUL-2004	31.318	-81.318	1	2.1	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0022	13-JUL-2004	31.292	-81.355	1	0.9	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0023	13-JUL-2004	31.276	-81.309	1	8.2	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0024	22-JUN-2004	31.227	-81.697	1	8.4	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0025	22-JUN-2004	31.2	-81.764	1	1.2	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0026	01-JUL-2004	31.107	-81.635	1	1.5	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0027	22-JUN-2004	31.077	-81.706	1	1.8	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0028	01-JUL-2004	31.053	-81.503	1	3.3	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0029	22-JUN-2004	31.064	-81.748	1	2.3	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0030	23-JUN-2004	31.018	-81.441	1	6.7	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0031	20-JUL-2004	30.738	-81.535	1	0.9	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0032	15-JUL-2004	30.722	-81.559	1	2.1	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0033	05-AUG-2004	31.958	-81.169	1	1.7	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0034	11-AUG-2004	31.922	-81.09	1	6.2	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0035	10-AUG-2004	31.857	-81.024	1	5.5	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0036	05-AUG-2004	31.858	-81.07	1	5.6	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0037	10-AUG-2004	31.852	-81.004	1	4.6	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0038	27-JUL-2004	31.702	-81.326	1	2.0	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0039	27-JUL-2004	31.592	-81.174	1	3.8	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0040	27-JUL-2004	31.59	-81.188	1	2.8	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0041	22-JUL-2004	31.541	-81.208	1	7.3	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0042	22-JUL-2004	31.54	-81.252	1	7.3	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0043	21-JUN-2004	31.095	-81.465	1	2.0	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0044	24-JUN-2004	30.975	-81.51	1	2.5	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0045	30-JUN-2004	30.97	-81.568	1	4.9	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0046	24-JUN-2004	30.987	-81.49	1	6.1	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0047	24-JUN-2004	30.934	-81.438	1	0.9	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0048	14-JUL-2004	30.842	-81.554	1	0.9	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0049	14-JUL-2004	30.738	-81.485	1	5.2	m	
National Coastal Assessment-Southeast/Georgia Dept. of Natural Resources-Coastal Resources	2004	GA04-0050	20-JUL-2004	30.709	-81.47	1	11.6	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0500	23-AUG-1997	36.518	-75.98	1	1.2	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0501	21-AUG-1997	36.461	-76.996	1	9.3	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0502	23-AUG-1997	36.413	-75.9	1	1.0	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0503	21-AUG-1997	36.396	-76.92	1	6.8	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0504	21-AUG-1997	36.375	-76.846	1	6.4	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0505	21-AUG-1997	36.363	-76.79	1	2.0	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0506	21-AUG-1997	36.292	-76.698	1	3.7	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0507	22-AUG-1997	36.235	-75.934	1	3.7	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0508	23-AUG-1997	36.23	-75.816	1	1.2	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0509	21-AUG-1997	36.218	-76.718	1	7.0	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0510	21-AUG-1997	36.174	-76.745	1	4.5	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0511	22-AUG-1997	36.149	-75.781	1	2.3	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0512	20-AUG-1997	36.137	-76.131	1	1.0	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0513	21-AUG-1997	36.117	-76.737	1	6.1	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0514	21-AUG-1997	36.083	-76.718	1	5.4	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0515	22-AUG-1997	36.087	-75.964	1	5.3	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0516	20-AUG-1997	36.072	-76.275	1	5.1	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0517	21-AUG-1997	36.026	-76.666	1	4.0	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0518	22-AUG-1997	35.952	-76.714	1	1.7	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0519	21-AUG-1997	35.917	-76.721	1	4.6	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0520	08-JUL-1997	35.92	-75.982	1	3.6	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0521	09-JUL-1997	35.824	-75.677	1	4.4	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0522	09-JUL-1997	35.739	-75.636	1	3.4	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0523	09-JUL-1997	35.698	-75.757	1	1.2	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0524	16-JUL-1997	35.5	-77.03	1	1.4	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0525	19-AUG-1997	35.448	-75.587	1	5.1	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0526	11-JUL-1997	35.429	-76.532	1	2.1	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0527	15-JUL-1997	35.406	-76.752	1	4.6	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0528	19-AUG-1997	35.412	-75.779	1	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0529	10-JUL-1997	35.406	-75.967	1	4.4	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0530	11-JUL-1997	35.388	-76.46	1	2.7	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0531	11-JUL-1997	35.376	-76.65	1	4.6	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0532	10-JUL-1997	35.359	-76.131	1	0.7	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0533	19-AUG-1997	35.37	-75.583	1	4.0	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0534	10-JUL-1997	35.339	-76.288	1	2.0	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0535	11-JUL-1997	35.321	-76.558	1	1.5	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0536	18-AUG-1997	35.322	-76.055	1	3.4	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0537	19-AUG-1997	35.275	-75.88	1	5.3	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0538	23-JUL-1997	35.237	-76.514	1	0.8	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0539	19-AUG-1997	35.236	-76.148	1	5.4	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0540	18-AUG-1997	35.233	-75.849	1	4.3	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0541	19-AUG-1997	35.192	-75.765	1	3.6	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0542	18-JUL-1997	35.071	-77.076	1	2.0	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0543	17-JUL-1997	35.089	-76.514	1	6.6	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0544	18-AUG-1997	35.077	-76.014	1	0.9	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0545	17-JUL-1997	35.0	-76.684	1	5.6	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0546	23-JUL-1997	34.975	-76.278	1	2.5	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0547	17-JUL-1997	34.967	-76.583	1	2.9	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1998	MA98-1041	16-JUL-1998	35.257	-77.29	1	0.8	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1998	MA98-1042	16-JUL-1998	35.229	-77.165	1	3.5	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1998	MA98-1043	16-JUL-1998	35.215	-77.133	1	2.0	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1998	MA98-1044	16-JUL-1998	35.204	-77.117	1	1.0	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1998	MA98-1045	16-JUL-1998	35.179	-77.092	1	1.9	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1998	MA98-1046	16-JUL-1998	35.162	-77.078	1	3.2	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1998	MA98-1047	15-JUL-1998	35.097	-77.029	1	2.9	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1998	MA98-1048	15-JUL-1998	35.07	-76.988	1	1.0	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1998	MA98-1049	15-JUL-1998	35.01	-76.941	1	3.0	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1998	MA98-1050	15-JUL-1998	35.003	-76.966	1	2.8	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1998	MA98-1051	15-JUL-1998	34.87	-76.897	1	3.9	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1998	MA98-1052	14-JUL-1998	34.988	-76.851	1	4.0	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1998	MA98-1053	14-JUL-1998	34.975	-76.775	1	1.2	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1998	MA98-1054	14-JUL-1998	34.947	-76.821	1	2.5	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1998	MA98-1055	14-JUL-1998	34.943	-76.772	1	3.0	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1998	MA98-1056	14-JUL-1998	34.995	-76.695	1	5.3	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1998	MA98-1057	13-JUL-1998	35.026	-76.601	1	5.9	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1998	MA98-1058	13-JUL-1998	35.103	-76.561	1	1.2	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1998	MA98-1059	13-JUL-1998	35.05	-76.502	1	6.5	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1998	MA98-1060	14-JUL-1998	35.011	-76.571	1	2.1	m	
National Coastal Assessment-Southeast/Environmental Protection Agency-Gulf Ecology Division	2000	NC00-0001	27-JUL-2000	36.442	-75.967	1	1.8	m	
National Coastal Assessment-Southeast/Environmental Protection Agency-Gulf Ecology Division	2000	NC00-0002	28-JUL-2000	36.115	-76.322	1	3.7	m	
National Coastal Assessment-Southeast/Environmental Protection Agency-Gulf Ecology Division	2000	NC00-0003	28-JUL-2000	35.964	-76.301	1	1.2	m	
National Coastal Assessment-Southeast/Environmental Protection Agency-Gulf Ecology Division	2000	NC00-0004	29-JUL-2000	35.953	-76.054	1	1.5	m	
National Coastal Assessment-Southeast/National Oceanic and Atmospheric Administration	2000	NC00-0005	17-AUG-2000	35.333	-76.176	1	1.0	m	
National Coastal Assessment-Southeast/National Oceanic and Atmospheric Administration	2000	NC00-0006	22-AUG-2000	34.982	-76.377	1	0.4	m	
National Coastal Assessment-Southeast/National Oceanic and Atmospheric Administration	2000	NC00-0007	22-AUG-2000	34.964	-76.454	1	0.5	m	
National Coastal Assessment-Southeast/National Oceanic and Atmospheric Administration	2000	NC00-0008	14-AUG-2000	34.889	-76.862	1	0.5	m	
National Coastal Assessment-Southeast/National Oceanic and Atmospheric Administration	2000	NC00-0009	21-AUG-2000	34.729	-77.104	1	0.3	m	
National Coastal Assessment-Southeast/National Oceanic and Atmospheric Administration	2000	NC00-0010	21-AUG-2000	34.627	-77.366	1	0.9	m	
National Coastal Assessment-Southeast/Environmental Protection Agency-Gulf Ecology Division	2000	NC00-0011	29-JUL-2000	35.96	-75.95	1	1.5	m	
National Coastal Assessment-Southeast/Environmental Protection Agency-Gulf Ecology Division	2000	NC00-0012	29-JUL-2000	35.768	-76.004	1	3.5	m	
National Coastal Assessment-Southeast/National Oceanic and Atmospheric Administration	2000	NC00-0013	16-AUG-2000	35.37	-76.603	1	1.6	m	
National Coastal Assessment-Southeast/National Oceanic and Atmospheric Administration	2000	NC00-0014	16-AUG-2000	35.301	-76.432	1	1.7	m	
National Coastal Assessment-Southeast/National Oceanic and Atmospheric Administration	2000	NC00-0015	16-AUG-2000	35.343	-76.59	1	1.4	m	
National Coastal Assessment-Southeast/National Oceanic and Atmospheric Administration	2000	NC00-0016	14-AUG-2000	35.021	-76.542	1	1.9	m	
National Coastal Assessment-Southeast/National Oceanic and Atmospheric Administration	2000	NC00-0017	16-AUG-2000	35.018	-76.619	1	1.7	m	
National Coastal Assessment-Southeast/National Oceanic and Atmospheric Administration	2000	NC00-0018	22-AUG-2000	34.939	-76.238	1	0.4	m	
National Coastal Assessment-Southeast/National Oceanic and Atmospheric Administration	2000	NC00-0019	18-AUG-2000	34.939	-76.75	1	1.4	m	
National Coastal Assessment-Southeast/National Oceanic and Atmospheric Administration	2000	NC00-0020	19-AUG-2000	34.775	-76.428	1	0.3	m	
National Coastal Assessment-Southeast/Environmental Protection Agency-Gulf Ecology Division	2000	NC00-0022	26-JUL-2000	36.085	-75.939	1	5.6	m	
National Coastal Assessment-Southeast/Environmental Protection Agency-Gulf Ecology Division	2000	NC00-0023	26-JUL-2000	36.071	-76.086	1	5.7	m	
National Coastal Assessment-Southeast/Environmental Protection Agency-Gulf Ecology Division	2000	NC00-0024	28-JUL-2000	36.01	-76.314	1	6.2	m	
National Coastal Assessment-Southeast/Environmental Protection Agency-Gulf Ecology Division	2000	NC00-0025	27-JUL-2000	35.988	-76.671	1	3.7	m	
National Coastal Assessment-Southeast/Environmental Protection Agency-Gulf Ecology Division	2000	NC00-0026	30-JUL-2000	35.629	-75.641	1	4.0	m	
National Coastal Assessment-Southeast/Environmental Protection Agency-Gulf Ecology Division	2000	NC00-0027	30-JUL-2000	35.499	-75.553	1	3.8	m	
National Coastal Assessment-Southeast/National Oceanic and Atmospheric Administration	2000	NC00-0028	17-AUG-2000	35.431	-75.834	1	1.9	m	
National Coastal Assessment-Southeast/National Oceanic and Atmospheric Administration	2000	NC00-0029	17-AUG-2000	35.361	-75.997	1	1.6	m	
National Coastal Assessment-Southeast/Environmental Protection Agency-Gulf Ecology Division	2000	NC00-0030	31-JUL-2000	35.22	-75.66	1	0.9	m	
National Coastal Assessment-Southeast/National Oceanic and Atmospheric Administration	2000	NC00-0031	17-AUG-2000	35.306	-76.223	1	1.3	m	
National Coastal Assessment-Southeast/National Oceanic and Atmospheric Administration	2000	NC00-0032	15-AUG-2000	35.169	-75.899	1	1.2	m	
National Coastal Assessment-Southeast/National Oceanic and Atmospheric Administration	2000	NC00-0033	15-AUG-2000	35.165	-76.226	1	1.9	m	
National Coastal Assessment-Southeast/National Oceanic and Atmospheric Administration	2000	NC00-0034	15-AUG-2000	35.136	-76.276	1	1.9	m	
National Coastal Assessment-Southeast/National Oceanic and Atmospheric Administration	2000	NC00-0035	15-AUG-2000	35.046	-76.161	1	1.0	m	
National Coastal Assessment-Southeast/USEPA, Science and Ecosystems Support Division	2001	NC01-0001	01-AUG-2001	36.432	-75.968	1	0.6	m	
National Coastal Assessment-Southeast/USEPA, Science and Ecosystems Support Division	2001	NC01-0002	02-AUG-2001	36.13	-76.346	1	1.1	m	
National Coastal Assessment-Southeast/USEPA, Science and Ecosystems Support Division	2001	NC01-0003	03-AUG-2001	35.935	-76.286	1	1.2	m	
National Coastal Assessment-Southeast/USEPA, Science and Ecosystems Support Division	2001	NC01-0004	05-AUG-2001	35.916	-76.061	1	1.2	m	
National Coastal Assessment-Southeast/USEPA, Science and Ecosystems Support Division	2001	NC01-0005	06-AUG-2001	35.339	-76.165	1	2.3	m	
National Coastal Assessment-Southeast/USEPA, Science and Ecosystems Support Division	2001	NC01-0006	05-AUG-2001	34.968	-76.341	1	1.4	m	
National Coastal Assessment-Southeast/USEPA, Science and Ecosystems Support Division	2001	NC01-0007	04-AUG-2001	34.926	-76.595	1	1.2	m	
National Coastal Assessment-Southeast/USEPA, Science and Ecosystems Support Division	2001	NC01-0008	03-AUG-2001	34.946	-76.915	1	1.0	m	
National Coastal Assessment-Southeast/USEPA, Science and Ecosystems Support Division	2001	NC01-0009	06-AUG-2001	34.693	-77.093	1	0.6	m	
National Coastal Assessment-Southeast/USEPA, Science and Ecosystems Support Division	2001	NC01-0010	07-AUG-2001	34.591	-77.418	1	1.8	m	
National Coastal Assessment-Southeast/USEPA, Science and Ecosystems Support Division	2001	NC01-0011	05-AUG-2001	35.982	-75.996	1	4.6	m	
National Coastal Assessment-Southeast/USEPA, Science and Ecosystems Support Division	2001	NC01-0012	05-AUG-2001	35.789	-76.03	1	3.2	m	
National Coastal Assessment-Southeast/USEPA, Science and Ecosystems Support Division	2001	NC01-0013	23-AUG-2001	35.363	-76.593	1	4.6	m	
National Coastal Assessment-Southeast/USEPA, Science and Ecosystems Support Division	2001	NC01-0014	31-JUL-2001	35.356	-76.387	1	1.7	m	
National Coastal Assessment-Southeast/USEPA, Science and Ecosystems Support Division	2001	NC01-0015	02-AUG-2001	35.339	-76.605	1	2.0	m	
National Coastal Assessment-Southeast/USEPA, Science and Ecosystems Support Division	2001	NC01-0016	24-AUG-2001	35.113	-76.54	1	4.6	m	
National Coastal Assessment-Southeast/USEPA, Science and Ecosystems Support Division	2001	NC01-0017	24-AUG-2001	34.98	-76.729	1	4.6	m	
National Coastal Assessment-Southeast/USEPA, Science and Ecosystems Support Division	2001	NC01-0018	05-AUG-2001	34.889	-76.322	1	1.6	m	
National Coastal Assessment-Southeast/USEPA, Science and Ecosystems Support Division	2001	NC01-0019	04-AUG-2001	34.941	-76.768	1	2.6	m	
National Coastal Assessment-Southeast/USEPA, Science and Ecosystems Support Division	2001	NC01-0020	08-AUG-2001	34.832	-76.361	1	0.9	m	
National Coastal Assessment-Southeast/USEPA, Science and Ecosystems Support Division	2001	NC01-0021	04-AUG-2001	36.267	-75.834	1	2.1	m	
National Coastal Assessment-Southeast/USEPA, Science and Ecosystems Support Division	2001	NC01-0022	04-AUG-2001	36.114	-75.927	1	4.9	m	
National Coastal Assessment-Southeast/USEPA, Science and Ecosystems Support Division	2001	NC01-0023	02-AUG-2001	36.072	-76.251	1	5.5	m	
National Coastal Assessment-Southeast/USEPA, Science and Ecosystems Support Division	2001	NC01-0025	31-JUL-2001	36.008	-76.556	1	2.7	m	
National Coastal Assessment-Southeast/USEPA, Science and Ecosystems Support Division	2001	NC01-0026	21-AUG-2001	35.611	-75.613	1	4.1	m	
National Coastal Assessment-Southeast/USEPA, Science and Ecosystems Support Division	2001	NC01-0027	08-AUG-2001	35.514	-75.695	1	5.5	m	
National Coastal Assessment-Southeast/USEPA, Science and Ecosystems Support Division	2001	NC01-0028	08-AUG-2001	35.437	-75.905	1	5.0	m	
National Coastal Assessment-Southeast/USEPA, Science and Ecosystems Support Division	2001	NC01-0029	07-AUG-2001	35.421	-76.001	1	2.7	m	
National Coastal Assessment-Southeast/USEPA, Science and Ecosystems Support Division	2001	NC01-0030	04-AUG-2001	35.271	-75.551	1	0.9	m	
National Coastal Assessment-Southeast/USEPA, Science and Ecosystems Support Division	2001	NC01-0031	23-AUG-2001	35.284	-76.334	1	1.8	m	
National Coastal Assessment-Southeast/USEPA, Science and Ecosystems Support Division	2001	NC01-0032	07-AUG-2001	35.256	-75.816	1	4.1	m	
National Coastal Assessment-Southeast/USEPA, Science and Ecosystems Support Division	2001	NC01-0033	23-AUG-2001	35.217	-76.203	1	4.3	m	
National Coastal Assessment-Southeast/USEPA, Science and Ecosystems Support Division	2001	NC01-0034	24-AUG-2001	35.058	-76.306	1	6.1	m	
National Coastal Assessment-Southeast/USEPA, Science and Ecosystems Support Division	2001	NC01-0035	07-AUG-2001	34.99	-76.167	1	0.5	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2002	NC02-0001	02-OCT-2002	36.396	-75.949	1	0.6	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2002	NC02-0002	19-SEP-2002	36.245	-76.131	1	2.5	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2002	NC02-0003	09-SEP-2002	36.299	-76.704	1	6.7	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2002	NC02-0004	19-SEP-2002	36.143	-75.984	1	4.0	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2002	NC02-0005	18-SEP-2002	36.123	-76.341	1	2.1	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2002	NC02-0006	18-SEP-2002	36.097	-76.196	1	1.2	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2002	NC02-0007	19-SEP-2002	35.971	-75.764	1	2.7	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2002	NC02-0008	18-SEP-2002	36.002	-76.232	1	5.5	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2002	NC02-0009	19-SEP-2002	35.88	-75.738	1	2.4	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2002	NC02-0010	23-SEP-2002	35.818	-75.58	1	0.8	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2002	NC02-0011	03-OCT-2002	35.746	-75.615	1	1.1	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2002	NC02-0012	09-SEP-2002	35.928	-76.717	1	3.0	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2002	NC02-0013	17-SEP-2002	35.789	-76.012	1	4.0	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2002	NC02-0014	24-SEP-2002	35.544	-75.476	1	0.6	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2002	NC02-0015	03-OCT-2002	35.578	-75.713	1	4.0	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2002	NC02-0016	04-NOV-2002	35.472	-75.892	1	4.9	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2002	NC02-0017	04-NOV-2002	35.408	-75.666	1	6.1	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2002	NC02-0018	05-SEP-2002	35.534	-76.506	1	2.7	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2002	NC02-0019	04-SEP-2002	35.435	-76.531	1	1.2	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2002	NC02-0020	08-NOV-2002	35.292	-75.705	1	3.0	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2002	NC02-0021	08-OCT-2002	35.335	-76.016	1	5.5	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2002	NC02-0022	08-NOV-2002	35.29	-75.828	1	4.0	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2002	NC02-0023	27-AUG-2002	35.475	-76.967	1	1.4	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2002	NC02-0024	03-SEP-2002	35.373	-76.377	1	2.4	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2002	NC02-0025	12-SEP-2002	35.331	-76.159	1	1.8	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2002	NC02-0026	29-AUG-2002	35.398	-76.726	1	4.7	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2002	NC02-0027	08-OCT-2002	35.239	-76.126	1	5.2	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2002	NC02-0028	03-OCT-2002	35.125	-76.296	1	6.1	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2002	NC02-0029	12-SEP-2002	35.159	-76.506	1	5.8	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2002	NC02-0030	03-OCT-2002	35.019	-76.428	1	1.9	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2002	NC02-0031	05-SEP-2002	34.949	-76.265	1	2.1	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2002	NC02-0032	29-AUG-2002	35.03	-76.953	1	2.6	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2002	NC02-0033	05-SEP-2002	34.869	-76.365	1	1.8	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2002	NC02-0034	04-SEP-2002	34.724	-76.696	1	2.7	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2002	NC02-0035	04-SEP-2002	34.712	-76.709	1	2.7	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2003	NC03-0001	26-AUG-2003	36.452	-76.011	1	0.7	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2003	NC03-0002	07-AUG-2003	36.201	-76.062	1	3.0	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2003	NC03-0003	15-AUG-2003	35.876	-75.621	1	0.9	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2003	NC03-0004	14-AUG-2003	35.858	-75.69	1	2.4	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2003	NC03-0005	08-JUL-2003	35.941	-76.644	1	2.1	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2003	NC03-0006	08-JUL-2003	35.919	-76.775	1	2.6	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2003	NC03-0007	30-JUL-2003	35.586	-75.814	1	1.5	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2003	NC03-0008	27-AUG-2003	35.009	-76.352	1	1.2	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2003	NC03-0009	16-JUL-2003	34.611	-77.365	1	0.2	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2003	NC03-0010	16-JUL-2003	34.143	-77.952	1	4.6	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2003	NC03-0011	12-AUG-2003	35.877	-76.027	1	3.0	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2003	NC03-0012	15-AUG-2003	35.811	-75.611	1	1.5	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2003	NC03-0013	29-JUL-2003	35.801	-76.004	1	3.4	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2003	NC03-0014	29-JUL-2003	35.691	-76.027	1	2.4	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2003	NC03-0015	21-AUG-2003	34.998	-76.271	1	0.1	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2003	NC03-0016	22-JUL-2003	35.006	-76.917	1	2.1	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2003	NC03-0017	08-AUG-2003	34.975	-76.733	1	4.9	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2003	NC03-0018	22-JUL-2003	34.979	-76.935	1	2.4	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2003	NC03-0019	09-JUL-2003	34.71	-76.483	1	0.9	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2003	NC03-0020	09-JUL-2003	34.704	-76.899	1	0.9	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2003	NC03-0021	26-AUG-2003	36.281	-75.817	1	0.6	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2003	NC03-0022	12-AUG-2003	36.092	-75.957	1	5.8	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2003	NC03-0023	05-AUG-2003	36.084	-76.14	1	5.8	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2003	NC03-0024	05-AUG-2003	36.026	-76.407	1	6.1	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2003	NC03-0025	14-AUG-2003	35.75	-75.622	1	1.8	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2003	NC03-0026	13-AUG-2003	35.541	-75.833	1	4.3	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2003	NC03-0027	17-JUL-2003	35.472	-75.969	1	3.7	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2003	NC03-0028	13-AUG-2003	35.462	-75.611	1	5.5	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2003	NC03-0029	20-AUG-2003	35.337	-75.778	1	5.3	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2003	NC03-0030	21-AUG-2003	35.313	-75.556	1	0.8	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2003	NC03-0031	15-JUL-2003	35.307	-76.196	1	3.4	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2003	NC03-0032	15-JUL-2003	35.291	-76.36	1	3.0	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2003	NC03-0033	20-AUG-2003	35.254	-75.902	1	5.6	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2003	NC03-0034	21-AUG-2003	35.072	-76.175	1	3.0	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2004	NC04-0001	15-SEP-2004	36.031	-76.125	1	4.9	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2004	NC04-0002	15-JUL-2004	35.064	-76.606	1	0.9	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2004	NC04-0003	08-JUL-2004	35.501	-76.62	1	0.7	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2004	NC04-0004	24-AUG-2004	36.096	-75.912	1	4.9	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2004	NC04-0005	05-AUG-2004	35.949	-75.988	1	4.0	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2004	NC04-0006	16-SEP-2004	36.138	-75.792	1	1.7	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2004	NC04-0007	07-JUL-2004	34.963	-76.806	1	3.0	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2004	NC04-0008	04-AUG-2004	36.081	-76.345	1	2.7	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2004	NC04-0009	01-SEP-2004	36.125	-76.099	1	3.4	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2004	NC04-0010	16-SEP-2004	36.038	-75.856	1	4.9	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2004	NC04-0011	17-AUG-2004	35.474	-75.579	1	5.2	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2004	NC04-0012	16-SEP-2004	35.08	-76.041	1	2.7	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2004	NC04-0013	15-JUL-2004	34.995	-76.655	1	3.0	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2004	NC04-0014	07-JUL-2004	34.717	-76.815	1	1.6	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2004	NC04-0015	22-SEP-2004	35.523	-75.763	1	5.2	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2004	NC04-0016	10-AUG-2004	35.36	-75.942	1	4.9	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2004	NC04-0017	12-JUL-2004	35.464	-76.509	1	1.2	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2004	NC04-0018	21-JUL-2004	35.262	-76.153	1	4.3	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2004	NC04-0019	30-JUL-2004	34.997	-76.513	1	0.7	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2004	NC04-0020	04-AUG-2004	36.042	-76.3	1	5.8	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2004	NC04-0021	17-AUG-2004	35.409	-75.586	1	4.9	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2004	NC04-0022	09-AUG-2004	35.138	-76.475	1	6.1	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2004	NC04-0023	11-AUG-2004	35.785	-75.572	1	1.1	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2004	NC04-0024	15-JUL-2004	35.665	-76.035	1	2.6	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2004	NC04-0025	05-AUG-2004	35.967	-75.851	1	1.7	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2004	NC04-0026	24-AUG-2004	36.161	-75.956	1	4.9	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2004	NC04-0027	19-AUG-2004	35.08	-76.421	1	0.5	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2004	NC04-0028	21-JUL-2004	35.312	-76.119	1	3.4	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2004	NC04-0029	05-AUG-2004	34.727	-77.36	1	1.2	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2004	NC04-0030	11-AUG-2004	35.656	-75.686	1	3.7	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2004	NC04-0031	23-SEP-2004	34.91	-76.261	1	0.6	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2004	NC04-0032	19-AUG-2004	35.067	-76.44	1	1.6	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2004	NC04-0033	10-AUG-2004	35.224	-75.975	1	6.4	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2004	NC04-0034	05-AUG-2004	34.155	-77.944	1	1.8	m	
National Coastal Assessment-Southeast/North Carolina Department of Natural Resources	2004	NC04-0035	30-JUL-2004	35.032	-76.398	1	3.7	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0001	08-AUG-2000	33.202	-79.187	1	4.5	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0002	11-JUL-2000	32.975	-79.911	1	11.3	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0003	27-JUN-2000	32.45	-80.503	1	5.0	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0004	20-JUN-2000	32.378	-80.706	1	1.9	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0005	20-JUN-2000	32.296	-80.648	1	6.4	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0006	08-AUG-2000	33.369	-79.248	1	2.4	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0007	18-JUL-2000	33.07	-79.474	1	2.3	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0008	28-JUN-2000	32.5	-80.445	1	5.5	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0009	28-JUN-2000	32.498	-80.516	1	8.3	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0010	01-AUG-2000	32.213	-80.878	1	4.0	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0011	08-AUG-2000	33.327	-79.279	1	2.9	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0012	08-AUG-2000	33.203	-79.272	1	3.2	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0013	26-JUL-2000	32.503	-80.358	1	8.8	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0014	28-JUN-2000	32.496	-80.576	1	4.8	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0015	21-JUN-2000	32.301	-80.802	1	10.6	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0016	19-JUL-2000	32.781	-79.877	1	1.2	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0017	09-AUG-2000	33.401	-79.24	1	4.7	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0018	25-JUL-2000	32.636	-80.269	1	6.1	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0019	05-JUL-2000	32.495	-80.8	1	6.7	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0020	21-JUN-2000	32.292	-80.726	1	2.0	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0021	12-JUL-2000	32.773	-80.075	1	3.0	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0022	15-AUG-2000	32.612	-80.478	1	7.3	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0023	21-JUN-2000	32.378	-80.791	1	8.9	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0024	20-JUN-2000	32.353	-80.653	1	6.3	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0025	21-JUN-2000	32.296	-80.759	1	4.5	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0026	09-AUG-2000	33.337	-79.176	1	4.1	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0027	11-JUL-2000	32.838	-79.947	1	6.6	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0028	15-AUG-2000	32.616	-80.166	1	5.0	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0029	05-JUL-2000	32.499	-80.825	1	5.6	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0030	01-AUG-2000	32.178	-80.772	1	4.0	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0031	02-AUG-2000	32.09	-80.915	1	3.1	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0032	26-JUL-2000	32.607	-80.537	1	4.4	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0033	25-JUL-2000	32.6	-80.203	1	2.0	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0034	27-JUN-2000	32.415	-80.598	1	1.4	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0035	18-JUL-2000	33.036	-79.395	1	3.2	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0036	20-JUN-2000	32.302	-80.584	1	1.6	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0037	25-JUL-2000	32.607	-80.274	1	1.5	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0038	05-JUL-2000	32.551	-80.834	1	2.4	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0039	19-JUL-2000	32.814	-79.755	1	2.9	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0040	18-JUL-2000	33.038	-79.492	1	3.0	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0041	26-JUL-2000	32.504	-80.306	1	1.3	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0042	19-JUL-2000	32.904	-79.626	1	2.4	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0043	12-JUL-2000	32.893	-80.108	1	1.9	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0044	28-JUN-2000	32.588	-80.449	1	1.0	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0045	19-JUL-2000	32.876	-79.696	1	1.1	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0046	11-JUL-2000	32.899	-79.901	1	2.6	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0047	01-AUG-2000	32.158	-80.843	1	4.3	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0048	12-JUL-2000	32.647	-80.058	1	0.6	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0049	27-JUN-2000	32.472	-80.508	1	1.8	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0050	12-JUL-2000	32.647	-79.988	1	3.0	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0051	16-AUG-2000	33.844	-78.607	1	2.0	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0052	01-AUG-2000	32.181	-80.822	1	3.1	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0053	25-JUL-2000	32.583	-80.187	1	1.7	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0054	27-JUN-2000	32.433	-80.601	1	1.0	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0055	11-JUL-2000	32.865	-79.922	1	1.0	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0056	16-AUG-2000	33.546	-79.021	1	2.1	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0057	02-AUG-2000	32.156	-80.952	1	2.6	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0058	02-AUG-2000	32.312	-80.917	1	1.8	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0059	05-JUL-2000	32.506	-80.758	1	1.3	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2000	SC00-0060	18-JUL-2000	33.047	-79.535	1	2.7	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0001	17-JUL-2001	33.27	-79.241	1	1.8	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0002	27-JUN-2001	32.924	-79.93	1	4.3	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0003	21-AUG-2001	32.449	-80.431	1	4.2	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0004	14-AUG-2001	32.405	-80.789	1	6.9	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0005	11-JUL-2001	32.231	-80.789	1	4.8	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0006	17-JUL-2001	33.291	-79.266	1	6.9	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0007	25-JUL-2001	32.919	-79.735	1	0.9	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0008	21-AUG-2001	32.451	-80.473	1	8.7	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0009	21-AUG-2001	32.534	-80.581	1	4.2	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0010	11-JUL-2001	32.244	-80.778	1	2.3	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0011	17-JUL-2001	33.333	-79.287	1	1.5	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0012	24-JUL-2001	33.176	-79.284	1	1.6	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0013	14-AUG-2001	32.5	-80.358	1	6.4	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0014	21-AUG-2001	32.489	-80.582	1	4.9	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0015	11-JUL-2001	32.309	-80.85	1	1.9	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0016	26-JUN-2001	32.757	-79.888	1	6.5	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0017	02-JUL-2001	33.872	-78.599	1	2.2	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0018	07-AUG-2001	32.637	-80.257	1	1.2	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0019	15-AUG-2001	32.521	-80.779	1	3.5	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0020	31-JUL-2001	32.303	-80.727	1	10.3	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0021	08-AUG-2001	32.677	-80.003	1	2.8	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0022	07-AUG-2001	32.596	-80.185	1	4.2	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0023	11-JUL-2001	32.359	-80.81	1	3.8	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0024	31-JUL-2001	32.387	-80.64	1	3.7	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0025	01-AUG-2001	32.397	-80.462	1	1.9	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0026	17-JUL-2001	33.314	-79.281	1	4.0	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0027	15-AUG-2001	32.871	-79.867	1	4.1	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0028	21-AUG-2001	32.447	-80.455	1	7.1	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0029	31-JUL-2001	32.456	-80.564	1	3.1	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0030	10-JUL-2001	32.165	-80.802	1	3.7	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0031	10-JUL-2001	32.217	-80.916	1	3.4	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0032	21-AUG-2001	32.592	-80.539	1	3.8	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0033	14-AUG-2001	32.434	-80.862	1	1.7	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0034	24-JUL-2001	33.04	-79.378	1	2.6	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0035	01-AUG-2001	32.313	-80.579	1	2.1	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0036	01-AUG-2001	32.317	-80.52	1	4.2	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0037	14-AUG-2001	32.513	-80.391	1	2.3	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0038	26-JUN-2001	32.89	-80.098	1	2.2	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0039	27-JUN-2001	32.898	-79.935	1	4.7	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0040	08-AUG-2001	32.621	-80.001	1	1.9	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0041	21-AUG-2001	32.521	-80.578	1	5.3	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0042	26-JUN-2001	32.716	-79.939	1	1.5	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0043	18-JUL-2001	33.349	-79.176	1	3.6	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0044	10-JUL-2001	32.162	-80.867	1	2.5	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0045	08-AUG-2001	32.633	-80.085	1	1.2	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0046	21-AUG-2001	32.489	-80.529	1	3.5	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0047	08-AUG-2001	32.66	-79.977	1	4.1	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0048	02-JUL-2001	33.857	-78.575	1	1.4	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0049	07-AUG-2001	32.565	-80.225	1	3.1	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0050	31-JUL-2001	32.42	-80.572	1	2.2	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0051	24-JUL-2001	33.192	-79.33	1	2.2	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0052	18-JUL-2001	33.532	-79.053	1	1.2	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0053	01-AUG-2001	32.325	-80.487	1	3.5	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0054	07-AUG-2001	32.645	-80.339	1	1.1	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2001	SC01-0055	25-JUL-2001	32.961	-79.615	1	2.1	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0001	18-JUN-2002	32.501	-80.502	1	16.7	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0002	07-AUG-2002	32.205	-80.801	1	2.6	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0003	09-JUL-2002	32.412	-80.682	1	5.6	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0004	16-JUL-2002	33.124	-79.269	1	1.4	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0005	18-JUN-2002	32.506	-80.556	1	7.6	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0006	21-AUG-2002	32.338	-80.475	1	5.0	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0007	19-JUN-2002	32.502	-80.637	1	2.6	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0008	17-JUL-2002	33.032	-79.473	1	3.1	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0009	06-AUG-2002	32.132	-80.829	1	14.8	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0010	17-JUL-2002	33.26	-79.258	1	3.5	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0011	06-AUG-2002	32.096	-80.948	1	6.2	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0012	17-JUL-2002	33.35	-79.276	1	4.4	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0013	25-JUN-2002	32.602	-80.242	1	3.5	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0014	13-AUG-2002	32.899	-79.842	1	6.9	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0015	31-JUL-2002	32.751	-79.895	1	0.9	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0016	09-JUL-2002	32.444	-80.805	1	3.9	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0017	23-JUL-2002	32.287	-80.712	1	10.8	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0018	20-AUG-2002	32.582	-80.621	1	6.5	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0019	07-AUG-2002	32.223	-80.784	1	4.4	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0020	23-JUL-2002	32.386	-80.84	1	2.7	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0021	09-JUL-2002	32.287	-80.655	1	10.0	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0022	23-JUL-2002	32.309	-80.804	1	6.7	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0023	16-JUL-2002	33.874	-78.586	1	2.8	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0024	26-JUN-2002	32.507	-80.457	1	2.2	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0025	31-JUL-2002	32.769	-79.874	1	5.9	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0026	26-JUN-2002	32.498	-80.444	1	4.1	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0027	13-AUG-2002	32.865	-79.961	1	12.5	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0028	26-JUN-2002	32.613	-80.404	1	2.8	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0029	31-JUL-2002	32.808	-79.965	1	2.3	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0030	10-JUL-2002	32.523	-80.844	1	2.1	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0032	21-AUG-2002	32.307	-80.548	1	4.1	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0033	14-AUG-2002	32.9	-79.635	1	2.0	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0034	25-JUN-2002	32.637	-80.362	1	4.3	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0035	31-JUL-2002	32.775	-79.824	1	2.3	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0036	10-JUL-2002	32.487	-80.804	1	1.8	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0037	30-JUL-2002	32.701	-79.915	1	1.8	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0038	10-JUL-2002	32.503	-80.846	1	2.2	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0039	09-JUL-2002	32.462	-80.665	1	1.2	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0040	19-JUN-2002	32.519	-80.586	1	2.2	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0041	17-JUL-2002	33.042	-79.393	1	2.6	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0042	19-JUN-2002	32.635	-80.587	1	2.0	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0043	26-JUN-2002	32.505	-80.377	1	3.1	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0044	25-JUN-2002	32.618	-80.332	1	2.1	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0045	06-AUG-2002	32.182	-80.754	1	1.8	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0046	18-JUN-2002	32.444	-80.597	1	2.7	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0047	13-AUG-2002	32.906	-79.93	1	5.1	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0048	14-AUG-2002	32.942	-79.788	1	1.4	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0049	06-AUG-2002	32.126	-81.004	1	3.8	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0050	23-JUL-2002	32.306	-80.928	1	1.3	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0051	30-JUL-2002	32.787	-80.081	1	1.8	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0052	30-JUL-2002	32.625	-80.025	1	3.0	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0053	21-AUG-2002	32.306	-80.557	1	4.0	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0054	18-JUN-2002	32.423	-80.603	1	3.7	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0055	07-AUG-2002	32.262	-80.796	1	2.8	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0056	13-AUG-2002	32.86	-79.851	1	2.4	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0057	14-AUG-2002	32.908	-79.64	1	1.7	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0058	10-JUL-2002	32.528	-80.794	1	1.8	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0059	19-JUN-2002	32.578	-80.514	1	2.2	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0060	30-JUL-2002	32.66	-79.966	1	3.0	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2002	SC02-0061	25-JUN-2002	32.577	-80.221	1	1.1	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0001	09-JUL-2003	32.526	-80.847	1	2.5	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0002	22-JUL-2003	32.317	-80.771	1	14.0	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0003	25-JUN-2003	32.379	-80.634	1	4.2	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0004	25-JUN-2003	32.286	-80.695	1	7.9	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0005	09-JUL-2003	32.494	-80.85	1	2.6	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0006	22-JUL-2003	32.297	-80.76	1	4.4	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0007	15-JUL-2003	32.54	-80.601	1	4.4	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0008	23-JUL-2003	32.154	-80.813	1	7.1	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0009	29-JUL-2003	32.681	-80.232	1	9.7	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0010	02-JUL-2003	32.991	-79.926	1	3.3	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0011	29-JUL-2003	32.676	-80.114	1	2.9	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0012	02-JUL-2003	32.926	-79.935	1	11.4	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0013	12-AUG-2003	32.561	-80.403	1	4.2	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0014	01-JUL-2003	32.784	-79.881	1	1.6	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0015	12-AUG-2003	32.772	-80.076	1	2.1	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0016	15-JUL-2003	32.474	-80.47	1	7.3	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0017	01-JUL-2003	32.759	-79.92	1	5.1	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0018	08-JUL-2003	32.645	-80.67	1	5.1	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0019	01-JUL-2003	32.791	-79.801	1	1.6	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0020	05-AUG-2003	33.29	-79.265	1	7.3	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0021	23-JUL-2003	32.142	-80.887	1	3.6	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0022	05-AUG-2003	33.341	-79.267	1	1.0	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0023	15-JUL-2003	32.519	-80.527	1	5.7	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0024	22-JUL-2003	32.176	-80.784	1	2.8	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0025	19-AUG-2003	32.364	-80.762	1	7.0	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0026	05-AUG-2003	33.145	-79.238	1	2.3	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0027	15-JUL-2003	32.486	-80.555	1	4.1	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0028	13-AUG-2003	33.532	-79.037	1	2.1	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0029	22-JUL-2003	32.327	-80.783	1	8.4	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0030	08-JUL-2003	32.598	-80.5	1	3.8	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0031	08-JUL-2003	32.617	-80.678	1	3.8	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0032	23-JUL-2003	32.115	-80.985	1	4.7	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0033	15-JUL-2003	32.439	-80.478	1	1.8	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0034	08-JUL-2003	32.553	-80.506	1	2.7	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0035	25-JUN-2003	32.421	-80.652	1	3.5	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0036	06-AUG-2003	33.047	-79.497	1	3.2	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0037	15-JUL-2003	32.506	-80.589	1	3.7	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0038	25-JUN-2003	32.395	-80.715	1	2.0	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0039	15-JUL-2003	32.433	-80.541	1	2.7	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0040	12-AUG-2003	32.897	-80.118	1	1.3	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0041	02-JUL-2003	32.988	-79.885	1	1.0	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0042	01-JUL-2003	32.72	-79.925	1	2.6	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0043	05-AUG-2003	33.199	-79.303	1	2.1	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0044	30-JUL-2003	32.617	-80.11	1	2.7	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0045	24-JUN-2003	32.334	-80.58	1	1.2	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0046	29-JUL-2003	32.699	-80.276	1	1.3	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0047	13-AUG-2003	32.829	-79.775	1	5.2	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0048	24-JUN-2003	32.371	-80.46	1	2.5	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0049	12-AUG-2003	32.546	-80.702	1	1.8	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0050	06-AUG-2003	33.06	-79.511	1	2.0	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0051	24-JUN-2003	32.29	-80.563	1	2.8	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0052	15-JUL-2003	32.487	-80.53	1	3.7	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0053	06-AUG-2003	33.088	-79.406	1	2.5	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0054	09-JUL-2003	32.425	-80.824	1	1.3	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0055	30-JUL-2003	32.699	-79.922	1	4.2	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0056	19-AUG-2003	32.222	-80.92	1	2.0	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0057	02-JUL-2003	32.827	-79.887	1	2.9	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0058	30-JUL-2003	32.616	-80.12	1	2.0	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0059	24-JUN-2003	32.342	-80.482	1	1.0	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2003	SC03-0060	06-AUG-2003	33.046	-79.483	1	1.3	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0001	29-JUN-2004	32.102	-81.007	1	9.9	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0002	03-AUG-2004	33.364	-79.268	1	2.7	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0003	30-JUN-2004	32.33	-80.721	1	5.4	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0004	03-AUG-2004	33.289	-79.281	1	3.6	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0005	28-JUL-2004	32.511	-80.361	1	6.2	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0006	10-AUG-2004	32.765	-79.907	1	4.6	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0007	17-AUG-2004	32.458	-80.445	1	8.7	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0008	11-AUG-2004	32.647	-80.013	1	1.6	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0009	17-AUG-2004	32.487	-80.481	1	10.6	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0010	08-JUL-2004	32.9	-79.955	1	5.1	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0011	17-AUG-2004	32.607	-80.484	1	6.3	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0012	10-AUG-2004	32.863	-79.719	1	2.5	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0013	13-JUL-2004	32.507	-80.595	1	1.8	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0014	20-JUL-2004	32.307	-80.61	1	3.7	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0015	21-JUL-2004	32.412	-80.794	1	10.0	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0016	03-AUG-2004	33.179	-79.26	1	3.6	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0017	14-JUL-2004	32.446	-80.533	1	3.1	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0018	18-AUG-2004	33.031	-79.418	1	2.7	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0019	13-JUL-2004	32.502	-80.655	1	3.3	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0020	29-JUN-2004	32.143	-80.832	1	2.5	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0021	27-JUL-2004	32.578	-80.203	1	9.6	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0022	04-AUG-2004	33.206	-79.19	1	3.6	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0023	27-JUL-2004	32.614	-80.259	1	6.9	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0024	08-JUL-2004	32.928	-79.793	1	2.3	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0025	21-JUL-2004	32.474	-80.836	1	5.0	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0026	30-JUN-2004	32.338	-80.752	1	8.2	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0027	13-JUL-2004	32.407	-80.67	1	5.6	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0028	29-JUN-2004	32.186	-80.733	1	2.6	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0029	21-JUL-2004	32.4	-80.813	1	5.2	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0030	30-JUN-2004	32.284	-80.742	1	10.3	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0031	21-JUL-2004	32.524	-80.819	1	3.1	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0032	18-AUG-2004	33.174	-79.379	1	2.6	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0033	29-JUN-2004	32.15	-80.967	1	3.3	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0034	04-AUG-2004	33.538	-79.039	1	1.6	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0035	14-JUL-2004	32.406	-80.604	1	2.3	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0036	03-AUG-2004	33.198	-79.313	1	2.9	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0037	13-JUL-2004	32.516	-80.727	1	3.5	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0038	08-JUL-2004	32.984	-79.907	1	2.5	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0039	07-JUL-2004	32.74	-79.9	1	1.6	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0040	11-AUG-2004	32.608	-80.126	1	1.5	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0041	20-JUL-2004	32.352	-80.501	1	2.0	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0042	27-JUL-2004	32.686	-80.217	1	2.8	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0043	10-AUG-2004	32.872	-79.692	1	3.1	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0044	27-JUL-2004	32.651	-80.209	1	2.2	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0045	10-AUG-2004	32.845	-79.754	1	3.5	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0046	17-AUG-2004	32.541	-80.509	1	4.1	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0047	20-JUL-2004	32.309	-80.537	1	1.3	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0048	17-AUG-2004	32.593	-80.67	1	5.9	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0049	18-AUG-2004	33.08	-79.428	1	2.0	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0050	14-JUL-2004	32.472	-80.618	1	1.2	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0051	18-AUG-2004	33.031	-79.583	1	2.8	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0052	20-JUL-2004	32.272	-80.627	1	1.6	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0053	28-JUL-2004	32.536	-80.335	1	2.8	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0054	30-JUN-2004	32.221	-80.822	1	1.5	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0055	28-JUL-2004	32.522	-80.311	1	2.1	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0056	28-JUL-2004	32.493	-80.325	1	2.2	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0057	14-JUL-2004	32.421	-80.601	1	2.9	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0058	11-AUG-2004	32.91	-80.138	1	1.0	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0059	07-JUL-2004	32.786	-80.129	1	5.2	m	
National Coastal Assessment-Southeast/South Carolina Department of Natural Resources	2004	SC04-0060	07-JUL-2004	32.734	-80.0	1	2.2	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0015	23-JUL-2001	36.548	-76.025	1	1.5	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0028	02-JUL-2002	36.55	-76.025	1	1.5	m	

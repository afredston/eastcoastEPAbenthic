
Search Parameters:Biogeographic Province in (Virginian))	
Data Group	Sampling Year	Station Name	Sampling Collection Date	Latitude Decimal Degrees	Longitude Decimal Degrees	Visit Number	Station Depth	Depth Units	
DE/MD Coastal Bays	1993	101	10-AUG-1993	38.588	-75.25	1	1.2	m	
DE/MD Coastal Bays	1993	102	10-AUG-1993	38.586	-75.273	1	0.9	m	
DE/MD Coastal Bays	1993	105	15-JUL-1993	38.584	-75.235	1	1.2	m	
DE/MD Coastal Bays	1993	105	30-SEP-1993	38.584	-75.235	2	1.2	m	
DE/MD Coastal Bays	1993	106	17-AUG-1993	38.593	-75.157	1	1.5	m	
DE/MD Coastal Bays	1993	107	04-AUG-1993	38.593	-75.17	1	1.2	m	
DE/MD Coastal Bays	1993	108	14-JUL-1993	38.593	-75.18	1	1.5	m	
DE/MD Coastal Bays	1993	108	24-SEP-1993	38.593	-75.18	2	1.5	m	
DE/MD Coastal Bays	1993	109	22-JUL-1993	38.591	-75.173	1	1.5	m	
DE/MD Coastal Bays	1993	109	24-SEP-1993	38.591	-75.173	2	1.5	m	
DE/MD Coastal Bays	1993	110	10-AUG-1993	38.588	-75.183	1	1.5	m	
DE/MD Coastal Bays	1993	111	24-AUG-1993	38.591	-75.154	1	1.8	m	
DE/MD Coastal Bays	1993	112	23-AUG-1993	38.588	-75.164	1	2.0	m	
DE/MD Coastal Bays	1993	113	26-AUG-1993	38.583	-75.16	1	1.2	m	
DE/MD Coastal Bays	1993	114	28-JUL-1993	38.582	-75.166	1	1.5	m	
DE/MD Coastal Bays	1993	115	28-JUL-1993	38.572	-75.192	1	1.8	m	
DE/MD Coastal Bays	1993	116	15-JUL-1993	38.588	-75.194	1	1.2	m	
DE/MD Coastal Bays	1993	116	24-SEP-1993	38.588	-75.194	2	1.2	m	
DE/MD Coastal Bays	1993	117	24-AUG-1993	38.588	-75.187	1	1.2	m	
DE/MD Coastal Bays	1993	118	17-AUG-1993	38.589	-75.204	1	0.8	m	
DE/MD Coastal Bays	1993	119	24-AUG-1993	38.583	-75.18	1	2.1	m	
DE/MD Coastal Bays	1993	120	26-AUG-1993	38.578	-75.176	1	1.2	m	
DE/MD Coastal Bays	1993	121	04-AUG-1993	38.575	-75.179	1	0.9	m	
DE/MD Coastal Bays	1993	122	10-AUG-1993	38.566	-75.204	1	1.8	m	
DE/MD Coastal Bays	1993	123	04-AUG-1993	38.592	-75.205	1	1.8	m	
DE/MD Coastal Bays	1993	124	10-AUG-1993	38.591	-75.216	1	1.5	m	
DE/MD Coastal Bays	1993	126	17-SEP-1993	38.591	-75.24	1	3.7	m	
DE/MD Coastal Bays	1993	127	21-SEP-1993	38.592	-75.186	1	0.9	m	
DE/MD Coastal Bays	1993	201	13-AUG-1993	38.37	-75.126	1	1.5	m	
DE/MD Coastal Bays	1993	202	26-JUL-1993	38.395	-75.129	1	1.5	m	
DE/MD Coastal Bays	1993	202	29-SEP-1993	38.395	-75.129	2	1.5	m	
DE/MD Coastal Bays	1993	203	16-JUL-1993	38.392	-75.124	1	1.5	m	
DE/MD Coastal Bays	1993	203	29-SEP-1993	38.392	-75.124	2	1.5	m	
DE/MD Coastal Bays	1993	204	13-AUG-1993	38.387	-75.119	1	1.5	m	
DE/MD Coastal Bays	1993	205	19-JUL-1993	38.388	-75.126	1	0.9	m	
DE/MD Coastal Bays	1993	205	29-SEP-1993	38.388	-75.126	2	0.9	m	
DE/MD Coastal Bays	1993	206	26-JUL-1993	38.383	-75.118	1	1.5	m	
DE/MD Coastal Bays	1993	206	29-SEP-1993	38.383	-75.118	2	1.5	m	
DE/MD Coastal Bays	1993	207	13-JUL-1993	38.378	-75.118	1	1.5	m	
DE/MD Coastal Bays	1993	207	29-SEP-1993	38.378	-75.118	2	1.5	m	
DE/MD Coastal Bays	1993	210	16-JUL-1993	38.379	-75.152	1	0.6	m	
DE/MD Coastal Bays	1993	211	13-AUG-1993	38.398	-75.117	1	1.5	m	
DE/MD Coastal Bays	1993	212	15-SEP-1993	38.398	-75.122	1	1.8	m	
DE/MD Coastal Bays	1993	213	27-AUG-1993	38.39	-75.117	1	1.5	m	
DE/MD Coastal Bays	1993	214	19-JUL-1993	38.387	-75.108	1	1.2	m	
DE/MD Coastal Bays	1993	214	29-SEP-1993	38.387	-75.108	2	1.2	m	
DE/MD Coastal Bays	1993	215	13-AUG-1993	38.404	-75.137	1	1.5	m	
DE/MD Coastal Bays	1993	216	23-JUL-1993	38.4	-75.134	1	1.2	m	
DE/MD Coastal Bays	1993	216	29-SEP-1993	38.4	-75.134	2	1.2	m	
DE/MD Coastal Bays	1993	217	23-JUL-1993	38.407	-75.146	1	1.2	m	
DE/MD Coastal Bays	1993	217	29-SEP-1993	38.407	-75.146	2	1.2	m	
DE/MD Coastal Bays	1993	218	16-JUL-1993	38.401	-75.141	1	0.9	m	
DE/MD Coastal Bays	1993	218	29-SEP-1993	38.401	-75.141	2	0.9	m	
DE/MD Coastal Bays	1993	219	13-AUG-1993	38.408	-75.153	1	1.2	m	
DE/MD Coastal Bays	1993	221	27-AUG-1993	38.412	-75.168	1	1.2	m	
DE/MD Coastal Bays	1993	223	19-JUL-1993	38.407	-75.179	1	1.2	m	
DE/MD Coastal Bays	1993	223	29-SEP-1993	38.407	-75.179	2	1.2	m	
DE/MD Coastal Bays	1993	224	31-AUG-1993	38.405	-75.176	1	0.9	m	
DE/MD Coastal Bays	1993	226	31-AUG-1993	38.383	-75.127	1	1.8	m	
DE/MD Coastal Bays	1993	227	31-AUG-1993	38.387	-75.115	1	1.5	m	
DE/MD Coastal Bays	1993	228	15-SEP-1993	38.398	-75.138	1	1.1	m	
DE/MD Coastal Bays	1993	301	07-SEP-1993	38.272	-75.177	1	0.9	m	
DE/MD Coastal Bays	1993	303	27-JUL-1993	38.232	-75.216	1	1.8	m	
DE/MD Coastal Bays	1993	304	22-SEP-1993	38.232	-75.228	1	1.8	m	
DE/MD Coastal Bays	1993	305	14-SEP-1993	38.237	-75.206	1	1.2	m	
DE/MD Coastal Bays	1993	306	12-AUG-1993	38.239	-75.217	1	1.5	m	
DE/MD Coastal Bays	1993	307	14-SEP-1993	38.226	-75.199	1	0.9	m	
DE/MD Coastal Bays	1993	308	14-SEP-1993	38.223	-75.209	1	1.8	m	
DE/MD Coastal Bays	1993	309	22-AUG-1993	38.226	-75.225	1	1.8	m	
DE/MD Coastal Bays	1993	310	28-AUG-1993	38.221	-75.22	1	2.1	m	
DE/MD Coastal Bays	1993	311	22-SEP-1993	38.219	-75.233	1	1.8	m	
DE/MD Coastal Bays	1993	312	14-SEP-1993	38.229	-75.231	1	1.8	m	
DE/MD Coastal Bays	1993	313	18-AUG-1993	38.262	-75.186	1	1.5	m	
DE/MD Coastal Bays	1993	314	27-JUL-1993	38.252	-75.198	1	1.2	m	
DE/MD Coastal Bays	1993	315	18-AUG-1993	38.279	-75.218	1	0.8	m	
DE/MD Coastal Bays	1993	316	18-AUG-1993	38.249	-75.184	1	1.5	m	
DE/MD Coastal Bays	1993	317	28-AUG-1993	38.232	-75.201	1	1.8	m	
DE/MD Coastal Bays	1993	318	20-AUG-1993	38.22	-75.208	1	2.1	m	
DE/MD Coastal Bays	1993	319	28-AUG-1993	38.215	-75.204	1	1.5	m	
DE/MD Coastal Bays	1993	320	22-AUG-1993	38.213	-75.211	1	1.5	m	
DE/MD Coastal Bays	1993	321	22-AUG-1993	38.207	-75.237	1	1.8	m	
DE/MD Coastal Bays	1993	322	22-AUG-1993	38.219	-75.235	1	1.5	m	
DE/MD Coastal Bays	1993	323	14-SEP-1993	38.215	-75.235	1	1.8	m	
DE/MD Coastal Bays	1993	324	27-JUL-1993	38.214	-75.245	1	1.5	m	
DE/MD Coastal Bays	1993	325	28-AUG-1993	38.21	-75.227	1	1.8	m	
DE/MD Coastal Bays	1993	401	21-SEP-1993	38.584	-75.068	1	1.5	m	
DE/MD Coastal Bays	1993	402	21-SEP-1993	38.578	-75.07	1	1.2	m	
DE/MD Coastal Bays	1993	403	03-SEP-1993	38.503	-75.067	1	1.2	m	
DE/MD Coastal Bays	1993	404	03-SEP-1993	38.502	-75.071	1	0.6	m	
DE/MD Coastal Bays	1993	405	09-SEP-1993	38.501	-75.087	1	0.8	m	
DE/MD Coastal Bays	1993	406	17-AUG-1993	38.642	-75.082	1	0.9	m	
DE/MD Coastal Bays	1993	407	15-JUL-1993	38.633	-75.087	1	0.6	m	
DE/MD Coastal Bays	1993	408	17-AUG-1993	38.638	-75.104	1	0.9	m	
DE/MD Coastal Bays	1993	409	04-AUG-1993	38.623	-75.089	1	3.4	m	
DE/MD Coastal Bays	1993	410	10-SEP-1993	38.672	-75.092	1	1.8	m	
DE/MD Coastal Bays	1993	411	21-AUG-1993	38.661	-75.095	1	1.8	m	
DE/MD Coastal Bays	1993	412	16-SEP-1993	38.65	-75.079	1	0.8	m	
DE/MD Coastal Bays	1993	413	14-JUL-1993	38.653	-75.089	1	0.9	m	
DE/MD Coastal Bays	1993	413	30-SEP-1993	38.653	-75.089	2	0.9	m	
DE/MD Coastal Bays	1993	414	19-AUG-1993	38.668	-75.12	1	1.2	m	
DE/MD Coastal Bays	1993	415	10-SEP-1993	38.664	-75.118	1	1.2	m	
DE/MD Coastal Bays	1993	416	26-AUG-1993	38.665	-75.126	1	1.5	m	
DE/MD Coastal Bays	1993	417	21-JUL-1993	38.655	-75.108	1	1.2	m	
DE/MD Coastal Bays	1993	417	30-SEP-1993	38.655	-75.108	2	1.2	m	
DE/MD Coastal Bays	1993	418	21-JUL-1993	38.643	-75.104	1	1.2	m	
DE/MD Coastal Bays	1993	418	30-SEP-1993	38.643	-75.104	2	1.2	m	
DE/MD Coastal Bays	1993	419	14-JUL-1993	38.662	-75.121	1	0.9	m	
DE/MD Coastal Bays	1993	419	30-SEP-1993	38.662	-75.121	2	0.9	m	
DE/MD Coastal Bays	1993	423	13-JUL-1993	38.605	-75.117	1	1.8	m	
DE/MD Coastal Bays	1993	423	24-SEP-1993	38.605	-75.117	2	1.8	m	
DE/MD Coastal Bays	1993	424	14-JUL-1993	38.596	-75.101	1	1.2	m	
DE/MD Coastal Bays	1993	424	30-SEP-1993	38.596	-75.101	2	1.2	m	
DE/MD Coastal Bays	1993	425	26-AUG-1993	38.585	-75.099	1	1.2	m	
DE/MD Coastal Bays	1993	426	21-JUL-1993	38.637	-75.117	1	1.5	m	
DE/MD Coastal Bays	1993	426	30-SEP-1993	38.637	-75.117	2	1.5	m	
DE/MD Coastal Bays	1993	427	16-SEP-1993	38.636	-75.114	1	0.6	m	
DE/MD Coastal Bays	1993	428	04-AUG-1993	38.63	-75.107	1	0.9	m	
DE/MD Coastal Bays	1993	429	21-JUL-1993	38.614	-75.104	1	0.9	m	
DE/MD Coastal Bays	1993	429	30-SEP-1993	38.614	-75.104	2	0.9	m	
DE/MD Coastal Bays	1993	430	21-JUL-1993	38.62	-75.126	1	0.6	m	
DE/MD Coastal Bays	1993	430	30-SEP-1993	38.62	-75.126	2	0.6	m	
DE/MD Coastal Bays	1993	433	27-AUG-1993	38.467	-75.059	1	0.6	m	
DE/MD Coastal Bays	1993	434	27-AUG-1993	38.486	-75.104	1	0.8	m	
DE/MD Coastal Bays	1993	435	16-AUG-1993	38.456	-75.062	1	1.8	m	
DE/MD Coastal Bays	1993	436	15-SEP-1993	38.457	-75.079	1	0.6	m	
DE/MD Coastal Bays	1993	438	21-AUG-1993	38.682	-75.098	1	2.1	m	
DE/MD Coastal Bays	1993	439	21-AUG-1993	38.691	-75.106	1	0.9	m	
DE/MD Coastal Bays	1993	440	14-JUL-1993	38.676	-75.107	1	1.5	m	
DE/MD Coastal Bays	1993	440	30-SEP-1993	38.676	-75.107	2	1.5	m	
DE/MD Coastal Bays	1993	441	19-AUG-1993	38.688	-75.137	1	1.4	m	
DE/MD Coastal Bays	1993	442	19-AUG-1993	38.679	-75.127	1	1.8	m	
DE/MD Coastal Bays	1993	444	28-JUL-1993	38.644	-75.143	1	0.9	m	
DE/MD Coastal Bays	1993	446	22-JUL-1993	38.639	-75.17	1	1.2	m	
DE/MD Coastal Bays	1993	446	30-SEP-1993	38.639	-75.17	2	1.2	m	
DE/MD Coastal Bays	1993	447	16-SEP-1993	38.64	-75.16	1	0.8	m	
DE/MD Coastal Bays	1993	448	15-JUL-1993	38.603	-75.145	1	1.8	m	
DE/MD Coastal Bays	1993	448	24-SEP-1993	38.603	-75.145	2	1.8	m	
DE/MD Coastal Bays	1993	450	21-JUL-1993	38.597	-75.138	1	1.8	m	
DE/MD Coastal Bays	1993	450	24-SEP-1993	38.597	-75.138	2	1.8	m	
DE/MD Coastal Bays	1993	451	17-SEP-1993	38.608	-75.098	1	2.4	m	
DE/MD Coastal Bays	1993	452	23-SEP-1993	38.601	-75.089	1	0.9	m	
DE/MD Coastal Bays	1993	454	21-SEP-1993	38.66	-75.086	1	1.8	m	
DE/MD Coastal Bays	1993	455	23-SEP-1993	38.67	-75.086	1	1.8	m	
DE/MD Coastal Bays	1993	501	13-JUL-1993	38.367	-75.111	1	1.2	m	
DE/MD Coastal Bays	1993	501	29-SEP-1993	38.367	-75.111	2	1.2	m	
DE/MD Coastal Bays	1993	502	12-JUL-1993	38.358	-75.137	1	0.9	m	
DE/MD Coastal Bays	1993	502	29-SEP-1993	38.358	-75.137	2	0.9	m	
DE/MD Coastal Bays	1993	503	13-JUL-1993	38.405	-75.09	1	2.4	m	
DE/MD Coastal Bays	1993	503	29-SEP-1993	38.405	-75.09	2	2.4	m	
DE/MD Coastal Bays	1993	504	13-JUL-1993	38.384	-75.087	1	1.2	m	
DE/MD Coastal Bays	1993	504	29-SEP-1993	38.384	-75.087	2	1.2	m	
DE/MD Coastal Bays	1993	505	13-JUL-1993	38.441	-75.078	1	1.8	m	
DE/MD Coastal Bays	1993	505	29-SEP-1993	38.441	-75.078	2	1.8	m	
DE/MD Coastal Bays	1993	506	23-JUL-1993	38.447	-75.079	1	1.2	m	
DE/MD Coastal Bays	1993	506	29-SEP-1993	38.447	-75.079	2	1.2	m	
DE/MD Coastal Bays	1993	507	23-JUL-1993	38.431	-75.102	1	1.2	m	
DE/MD Coastal Bays	1993	507	29-SEP-1993	38.431	-75.102	2	1.2	m	
DE/MD Coastal Bays	1993	508	20-AUG-1993	38.3	-75.121	1	0.8	m	
DE/MD Coastal Bays	1993	509	20-AUG-1993	38.235	-75.158	1	1.2	m	
DE/MD Coastal Bays	1993	510	20-JUL-1993	38.154	-75.226	1	1.8	m	
DE/MD Coastal Bays	1993	510	28-SEP-1993	38.154	-75.226	2	1.8	m	
DE/MD Coastal Bays	1993	512	22-SEP-1993	38.142	-75.248	1	2.1	m	
DE/MD Coastal Bays	1993	513	20-JUL-1993	38.179	-75.251	1	1.8	m	
DE/MD Coastal Bays	1993	513	28-SEP-1993	38.179	-75.251	2	1.8	m	
DE/MD Coastal Bays	1993	514	27-JUL-1993	38.154	-75.261	1	1.5	m	
DE/MD Coastal Bays	1993	515	14-SEP-1993	38.177	-75.224	1	1.8	m	
DE/MD Coastal Bays	1993	516	20-JUL-1993	38.169	-75.216	1	1.2	m	
DE/MD Coastal Bays	1993	516	28-SEP-1993	38.169	-75.216	2	1.2	m	
DE/MD Coastal Bays	1993	517	22-SEP-1993	38.173	-75.229	1	1.8	m	
DE/MD Coastal Bays	1993	520	25-AUG-1993	38.086	-75.252	1	1.2	m	
DE/MD Coastal Bays	1993	521	20-JUL-1993	38.22	-75.171	1	1.5	m	
DE/MD Coastal Bays	1993	521	28-SEP-1993	38.22	-75.171	2	1.5	m	
DE/MD Coastal Bays	1993	522	27-JUL-1993	38.209	-75.184	1	1.8	m	
DE/MD Coastal Bays	1993	523	22-AUG-1993	38.191	-75.191	1	1.2	m	
DE/MD Coastal Bays	1993	524	20-AUG-1993	38.201	-75.224	1	1.8	m	
DE/MD Coastal Bays	1993	525	27-JUL-1993	38.183	-75.247	1	1.8	m	
DE/MD Coastal Bays	1993	526	28-AUG-1993	38.194	-75.164	1	0.6	m	
DE/MD Coastal Bays	1993	527	28-AUG-1993	38.179	-75.18	1	0.9	m	
DE/MD Coastal Bays	1993	530	20-JUL-1993	38.048	-75.265	1	1.5	m	
DE/MD Coastal Bays	1993	530	28-SEP-1993	38.048	-75.265	2	1.5	m	
DE/MD Coastal Bays	1993	531	20-SEP-1993	38.079	-75.261	1	1.5	m	
DE/MD Coastal Bays	1993	532	25-AUG-1993	38.068	-75.261	1	0.8	m	
DE/MD Coastal Bays	1993	533	05-AUG-1993	38.07	-75.284	1	1.8	m	
DE/MD Coastal Bays	1993	536	05-AUG-1993	38.109	-75.261	1	2.1	m	
DE/MD Coastal Bays	1993	537	13-SEP-1993	38.115	-75.274	1	2.1	m	
DE/MD Coastal Bays	1993	538	11-AUG-1993	38.05	-75.288	1	1.2	m	
DE/MD Coastal Bays	1993	540	25-AUG-1993	38.038	-75.304	1	2.1	m	
DE/MD Coastal Bays	1993	541	20-JUL-1993	38.117	-75.292	1	0.9	m	
DE/MD Coastal Bays	1993	541	28-SEP-1993	38.117	-75.292	2	0.9	m	
DE/MD Coastal Bays	1993	543	05-AUG-1993	38.084	-75.322	1	1.2	m	
DE/MD Coastal Bays	1993	545	05-AUG-1993	38.075	-75.34	1	0.9	m	
DE/MD Coastal Bays	1993	547	24-SEP-1993	38.032	-75.366	1	1.2	m	
DE/MD Coastal Bays	1993	548	24-SEP-1993	38.055	-75.329	1	0.9	m	
DE/MD Coastal Bays	1993	549	26-JUL-1993	38.415	-75.073	1	1.5	m	
DE/MD Coastal Bays	1993	549	29-SEP-1993	38.415	-75.073	2	1.5	m	
DE/MD Coastal Bays	1993	550	26-JUL-1993	38.414	-75.087	1	1.5	m	
DE/MD Coastal Bays	1993	550	29-SEP-1993	38.414	-75.087	2	1.5	m	
DE/MD Coastal Bays	1993	551	22-SEP-1993	38.139	-75.284	1	0.9	m	
DE/MD Coastal Bays	1993	552	24-SEP-1993	38.029	-75.322	1	1.8	m	
DE/MD Coastal Bays	1993	553	23-SEP-1993	38.432	-75.072	1	1.5	m	
DE/MD Coastal Bays	1993	554	22-SEP-1993	38.111	-75.257	1	2.1	m	
DE/MD Coastal Bays	1993	555	22-SEP-1993	38.106	-75.231	1	1.8	m	
DE/MD Coastal Bays	1993	601	21-SEP-1993	38.628	-75.127	1	1.8	m	
DE/MD Coastal Bays	1993	603	13-JUL-1993	38.437	-75.078	1	3.4	m	
DE/MD Coastal Bays	1993	603	29-SEP-1993	38.437	-75.078	2	3.4	m	
DE/MD Coastal Bays	1993	604	26-JUL-1993	38.428	-75.06	1	1.8	m	
DE/MD Coastal Bays	1993	604	29-SEP-1993	38.428	-75.06	2	1.8	m	
DE/MD Coastal Bays	1993	605	16-SEP-1993	38.639	-75.159	1	1.5	m	
DE/MD Coastal Bays	1993	606	21-SEP-1993	38.617	-75.144	1	1.8	m	
DE/MD Coastal Bays	1993	610	21-AUG-1993	38.701	-75.111	1	2.1	m	
DE/MD Coastal Bays	1993	611	27-JUL-1993	38.233	-75.181	1	1.2	m	
DE/MD Coastal Bays	1993	612	28-JUL-1993	38.605	-75.077	1	1.8	m	
DE/MD Coastal Bays	1993	613	31-AUG-1993	38.464	-75.097	1	1.2	m	
DE/MD Coastal Bays	1993	614	27-JUL-1993	38.295	-75.132	1	2.7	m	
DE/MD Coastal Bays	1993	615	31-AUG-1993	38.465	-75.085	1	1.8	m	
DE/MD Coastal Bays	1993	616	19-JUL-1993	38.418	-75.171	1	0.9	m	
DE/MD Coastal Bays	1993	616	29-SEP-1993	38.418	-75.171	2	0.9	m	
DE/MD Coastal Bays	1993	617	10-AUG-1993	38.576	-75.095	1	1.8	m	
DE/MD Coastal Bays	1993	618	19-AUG-1993	38.689	-75.122	1	2.7	m	
DE/MD Coastal Bays	1993	619	21-AUG-1993	38.697	-75.084	1	0.9	m	
DE/MD Coastal Bays	1993	620	16-JUL-1993	38.374	-75.135	1	1.5	m	
DE/MD Coastal Bays	1993	620	29-SEP-1993	38.374	-75.135	2	1.5	m	
DE/MD Coastal Bays	1993	621	21-SEP-1993	38.592	-75.065	1	0.9	m	
DE/MD Coastal Bays	1993	622	14-JUL-1993	38.628	-75.11	1	0.9	m	
DE/MD Coastal Bays	1993	622	24-SEP-1993	38.628	-75.11	2	0.9	m	
DE/MD Coastal Bays	1993	623	19-JUL-1993	38.355	-75.118	1	0.9	m	
DE/MD Coastal Bays	1993	623	29-SEP-1993	38.355	-75.118	2	0.9	m	
DE/MD Coastal Bays	1993	624	27-AUG-1993	38.454	-75.057	1	0.8	m	
DE/MD Coastal Bays	1993	625	04-AUG-1993	38.56	-75.092	1	0.9	m	
DE/MD Coastal Bays	1993	626	21-AUG-1993	38.697	-75.097	1	1.2	m	
DE/MD Coastal Bays	1993	627	21-AUG-1993	38.691	-75.134	1	1.5	m	
DE/MD Coastal Bays	1993	628	29-SEP-1993	38.389	-75.071	1	2.1	m	
DE/MD Coastal Bays	1993	701	22-JUL-1993	38.695	-75.096	1	1.8	m	
DE/MD Coastal Bays	1993	701	28-JUL-1993	38.695	-75.096	2	1.8	m	
DE/MD Coastal Bays	1993	701	19-AUG-1993	38.695	-75.096	3	0.9	m	
DE/MD Coastal Bays	1993	701	24-AUG-1993	38.695	-75.096	4	1.8	m	
DE/MD Coastal Bays	1993	702	19-AUG-1993	38.662	-75.076	1			
DE/MD Coastal Bays	1993	702	24-AUG-1993	38.662	-75.076	2	0.8	m	
DE/MD Coastal Bays	1993	702	10-SEP-1993	38.662	-75.076	3	0.6	m	
DE/MD Coastal Bays	1993	702	16-SEP-1993	38.662	-75.076	4	0.8	m	
DE/MD Coastal Bays	1993	703	04-AUG-1993	38.598	-75.117	1	2.1	m	
DE/MD Coastal Bays	1993	703	10-AUG-1993	38.598	-75.117	2	2.4	m	
DE/MD Coastal Bays	1993	703	26-AUG-1993	38.598	-75.117	3	2.1	m	
DE/MD Coastal Bays	1993	703	30-AUG-1993	38.598	-75.117	4	2.1	m	
DE/MD Coastal Bays	1993	704	15-JUL-1993	38.583	-75.217	1	1.8	m	
DE/MD Coastal Bays	1993	704	21-JUL-1993	38.583	-75.217	2	1.5	m	
DE/MD Coastal Bays	1993	704	17-AUG-1993	38.583	-75.217	3	1.5	m	
DE/MD Coastal Bays	1993	704	23-AUG-1993	38.583	-75.217	4	1.2	m	
DE/MD Coastal Bays	1993	704	24-SEP-1993	38.583	-75.217	2	1.8	m	
DE/MD Coastal Bays	1993	705	09-AUG-1993	38.517	-75.063	1	0.9	m	
DE/MD Coastal Bays	1993	705	16-AUG-1993	38.517	-75.063	2	1.5	m	
DE/MD Coastal Bays	1993	705	03-SEP-1993	38.517	-75.063	3	0.9	m	
DE/MD Coastal Bays	1993	705	09-SEP-1993	38.517	-75.063	4	1.1	m	
DE/MD Coastal Bays	1993	706	09-AUG-1993	38.414	-75.175	1	0.9	m	
DE/MD Coastal Bays	1993	706	16-AUG-1993	38.414	-75.175	2	1.2	m	
DE/MD Coastal Bays	1993	706	03-SEP-1993	38.414	-75.175	3	1.2	m	
DE/MD Coastal Bays	1993	706	09-SEP-1993	38.414	-75.175	4	1.1	m	
DE/MD Coastal Bays	1993	707	12-AUG-1993	38.298	-75.181	1	0.8	m	
DE/MD Coastal Bays	1993	707	18-AUG-1993	38.298	-75.181	2	0.8	m	
DE/MD Coastal Bays	1993	707	02-SEP-1993	38.298	-75.181	3	0.9	m	
DE/MD Coastal Bays	1993	707	07-SEP-1993	38.298	-75.181	4	0.9	m	
DE/MD Coastal Bays	1993	708	12-AUG-1993	38.126	-75.235	1	1.8	m	
DE/MD Coastal Bays	1993	708	18-AUG-1993	38.126	-75.235	2	2.1	m	
DE/MD Coastal Bays	1993	708	02-SEP-1993	38.126	-75.235	3	2.1	m	
DE/MD Coastal Bays	1993	708	07-SEP-1993	38.126	-75.235	4	2.4	m	
DE/MD Coastal Bays	1993	709	05-AUG-1993	38.083	-75.225	1	1.2	m	
DE/MD Coastal Bays	1993	709	12-AUG-1993	38.083	-75.225	2	1.2	m	
DE/MD Coastal Bays	1993	709	25-AUG-1993	38.083	-75.225	3	1.5	m	
DE/MD Coastal Bays	1993	709	30-AUG-1993	38.083	-75.225	4	1.8	m	
DE/MD Coastal Bays	1993	710	11-AUG-1993	38.02	-75.349	1	1.8	m	
DE/MD Coastal Bays	1993	710	18-AUG-1993	38.02	-75.349	2	2.1	m	
DE/MD Coastal Bays	1993	710	02-SEP-1993	38.02	-75.349	3	2.1	m	
DE/MD Coastal Bays	1993	710	07-SEP-1993	38.02	-75.349	4	2.1	m	
DE/MD Coastal Bays	1993	711	05-AUG-1993	38.063	-75.312	1	1.2	m	
DE/MD Coastal Bays	1993	711	13-SEP-1993	38.063	-75.312	2	1.7	m	
DE/MD Coastal Bays	1993	711	20-SEP-1993	38.063	-75.312	3			
DE/MD Coastal Bays	1993	711	24-SEP-1993	38.063	-75.312	4	1.8	m	
DE/MD Coastal Bays	1993	712	20-JUL-1993	38.088	-75.288	1	1.8	m	
DE/MD Coastal Bays	1993	712	13-SEP-1993	38.088	-75.288	2	1.8	m	
DE/MD Coastal Bays	1993	712	20-SEP-1993	38.088	-75.288	3	1.8	m	
DE/MD Coastal Bays	1993	712	24-SEP-1993	38.088	-75.288	4	1.5	m	
DE/MD Coastal Bays	1993	713	20-JUL-1993	38.04	-75.286	1	1.2	m	
DE/MD Coastal Bays	1993	713	25-AUG-1993	38.04	-75.286	2	1.8	m	
DE/MD Coastal Bays	1993	713	13-SEP-1993	38.04	-75.286	3	1.8	m	
DE/MD Coastal Bays	1993	713	20-SEP-1993	38.04	-75.286	4	1.8	m	
DE/MD Coastal Bays	1993	714	05-AUG-1993	38.132	-75.206	1	1.2	m	
DE/MD Coastal Bays	1993	714	25-AUG-1993	38.132	-75.206	2	1.2	m	
DE/MD Coastal Bays	1993	714	13-SEP-1993	38.132	-75.206	3	0.9	m	
DE/MD Coastal Bays	1993	714	20-SEP-1993	38.132	-75.206	4	1.5	m	
DE/MD Coastal Bays	1993	715	27-AUG-1993	38.407	-75.172	1	1.1	m	
DE/MD Coastal Bays	1993	715	31-AUG-1993	38.407	-75.172	2	0.9	m	
DE/MD Coastal Bays	1993	715	09-SEP-1993	38.407	-75.172	3	1.2	m	
DE/MD Coastal Bays	1993	715	15-SEP-1993	38.407	-75.172	4	1.1	m	
DE/MD Coastal Bays	1993	716	27-AUG-1993	38.486	-75.084	1	1.1	m	
DE/MD Coastal Bays	1993	716	31-AUG-1993	38.486	-75.084	2	0.9	m	
DE/MD Coastal Bays	1993	716	08-SEP-1993	38.486	-75.084	3	0.9	m	
DE/MD Coastal Bays	1993	716	15-SEP-1993	38.486	-75.084	4	1.1	m	
DE/MD Coastal Bays	1993	717	15-JUL-1993	38.617	-75.1	1	1.2	m	
DE/MD Coastal Bays	1993	717	21-JUL-1993	38.617	-75.1	2	0.9	m	
DE/MD Coastal Bays	1993	717	17-AUG-1993	38.617	-75.1	3	1.2	m	
DE/MD Coastal Bays	1993	717	23-AUG-1993	38.617	-75.1	4	1.2	m	
DE/MD Coastal Bays	1993	717	24-SEP-1993	38.617	-75.1	2	1.2	m	
DE/MD Coastal Bays	1993	718	04-AUG-1993	38.585	-75.265	1	1.2	m	
DE/MD Coastal Bays	1993	718	10-AUG-1993	38.585	-75.265	2	0.9	m	
DE/MD Coastal Bays	1993	718	24-AUG-1993	38.585	-75.265	3	0.9	m	
DE/MD Coastal Bays	1993	718	30-AUG-1993	38.585	-75.265	4	0.9	m	
DE/MD Coastal Bays	1993	719	22-JUL-1993	38.655	-75.177	1	0.9	m	
DE/MD Coastal Bays	1993	719	28-JUL-1993	38.655	-75.177	2	0.8	m	
DE/MD Coastal Bays	1993	719	19-AUG-1993	38.655	-75.177	3	0.9	m	
DE/MD Coastal Bays	1993	719	24-AUG-1993	38.655	-75.177	4			
DE/MD Coastal Bays	1993	720	17-AUG-1993	38.655	-75.125	1	1.2	m	
DE/MD Coastal Bays	1993	720	26-AUG-1993	38.655	-75.125	2	0.8	m	
DE/MD Coastal Bays	1993	720	10-SEP-1993	38.655	-75.125	3	0.9	m	
DE/MD Coastal Bays	1993	720	16-SEP-1993	38.655	-75.125	4	0.8	m	
R-EMAP Region 2 1993-94	1993	BA002	03-OCT-1993	40.562	-73.686	1	12.5	m	
R-EMAP Region 2 1993-94	1993	BA005	03-OCT-1993	40.513	-73.584	1	20.7	m	
R-EMAP Region 2 1993-94	1993	BA007	04-OCT-1993	40.482	-73.764	1	26.8	m	
R-EMAP Region 2 1993-94	1993	BA010	04-OCT-1993	40.469	-73.915	1	18.9	m	
R-EMAP Region 2 1993-94	1993	BA012	04-OCT-1993	40.435	-73.688	1	26.2	m	
R-EMAP Region 2 1993-94	1993	BA014	04-OCT-1993	40.413	-73.797	1	35.7	m	
R-EMAP Region 2 1993-94	1993	BA016	04-OCT-1993	40.398	-73.876	1	22.6	m	
R-EMAP Region 2 1993-94	1993	BA017	04-OCT-1993	40.384	-73.56	1	26.2	m	
R-EMAP Region 2 1993-94	1993	BA021	05-OCT-1993	40.33	-73.517	1	27.1	m	
R-EMAP Region 2 1993-94	1993	BA025	28-SEP-1993	40.301	-73.941	1	16.8	m	
R-EMAP Region 2 1993-94	1993	BA026	05-OCT-1993	40.275	-73.564	1	30.2	m	
R-EMAP Region 2 1993-94	1993	BA030	05-OCT-1993	40.219	-73.61	1	31.7	m	
R-EMAP Region 2 1993-94	1993	BA033	04-OCT-1993	40.193	-73.853	1	23.8	m	
R-EMAP Region 2 1993-94	1993	BA035	04-OCT-1993	40.177	-73.735	1	41.1	m	
R-EMAP Region 2 1993-94	1994	BA102	11-AUG-1994	40.562	-73.836	1	9.8	m	
R-EMAP Region 2 1993-94	1994	BA103	30-AUG-1994	40.541	-73.932	1	8.8	m	
R-EMAP Region 2 1993-94	1994	BA104	11-AUG-1994	40.499	-73.545	1	20.4	m	
R-EMAP Region 2 1993-94	1994	BA105	11-AUG-1994	40.486	-73.507	1	21.9	m	
R-EMAP Region 2 1993-94	1994	BA106	30-AUG-1994	40.473	-73.99	1	7.0	m	
R-EMAP Region 2 1993-94	1994	BA107	11-AUG-1994	40.386	-73.942	1	14.3	m	
R-EMAP Region 2 1993-94	1994	BA108	11-AUG-1994	40.381	-73.823	1	32.6	m	
R-EMAP Region 2 1993-94	1994	BA109	10-AUG-1994	40.336	-73.719	1	25.9	m	
R-EMAP Region 2 1993-94	1994	BA110	10-AUG-1994	40.307	-73.625	1	26.2	m	
R-EMAP Region 2 1993-94	1994	BA111	10-AUG-1994	40.302	-73.888	1	20.7	m	
R-EMAP Region 2 1993-94	1994	BA112	10-AUG-1994	40.298	-73.734	1	26.8	m	
R-EMAP Region 2 1993-94	1994	BA113	15-SEP-1994	40.251	-73.988	1	5.8	m	
R-EMAP Region 2 1993-94	1994	BA114	10-AUG-1994	40.188	-73.802	1	30.5	m	
R-EMAP Region 2 1993-94	1994	BA115	11-AUG-1994	40.575	-73.781	1	10.4	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	BU01-0001-A	22-AUG-2001	41.604	-70.643	1	2.9	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	BU01-0002-C	22-AUG-2001	41.757	-70.712	1	8.2	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	BU01-0007-A	07-AUG-2001	41.695	-70.751	1	3.1	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	BU01-0013-C	22-AUG-2001	41.566	-70.651	1	2.5	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	BU01-0015-A	21-AUG-2001	41.591	-70.956	1	1.0	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	BU01-0016-C	21-AUG-2001	41.557	-71.067	1	1.9	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	BU01-0018-A	08-AUG-2001	41.551	-70.838	1	10.0	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	BU01-0019-A	07-AUG-2001	41.52	-70.759	1	15.0	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	BU01-0020-A	07-AUG-2001	41.508	-70.732	1	13.1	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	BU01-0021-A	08-AUG-2001	41.509	-70.958	1	9.4	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	BU01-0026-B	08-AUG-2001	41.463	-71.0	1	21.2	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	BU01-0029-A	08-AUG-2001	41.474	-71.114	1	15.9	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	BU01-0030-A	08-AUG-2001	41.435	-70.972	1	19.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	CT00-0001-A	17-AUG-2000	41.151	-73.22	1	1.8	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	CT00-0003-A	04-AUG-2000	41.288	-73.071	1	8.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	CT00-0005-A	18-SEP-2000	41.274	-72.327	1	1.5	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	CT00-0007-A	10-AUG-2000	41.298	-73.066	1	10.6	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	CT00-0009-A	03-AUG-2000	41.292	-72.348	1	4.6	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	CT00-0009-A	29-AUG-2000	41.292	-72.348	2	5.1	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	CT00-0009-A	31-AUG-2000	41.292	-72.348	3	5.1	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	CT00-0011-B	01-SEP-2000	41.331	-72.086	1	6.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	CT00-0013-B	03-AUG-2000	41.403	-72.426	1	5.3	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	CT00-0013-B	29-AUG-2000	41.403	-72.426	2	2.8	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	CT00-0015-A	06-SEP-2000	41.336	-72.176	1	2.4	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	CT00-0017-A	05-SEP-2000	41.348	-71.97	1	1.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	CT00-0021-A	07-AUG-2000	40.963	-73.623	1	15.9	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	CT00-0023-A	08-AUG-2000	40.979	-73.56	1	24.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	CT00-0025-A	08-AUG-2000	41.009	-73.513	1	13.8	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	CT00-0029-A	16-AUG-2000	41.12	-73.162	1	10.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	CT00-0035-A	25-JUL-2000	41.209	-72.908	1	10.9	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	CT00-0037-A	25-JUL-2000	41.196	-72.775	1	14.5	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	CT00-0039-A	25-JUL-2000	41.242	-72.665	1	10.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	CT00-0041-A	25-JUL-2000	41.246	-72.468	1	15.4	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	CT00-0045-A	21-JUL-2000	41.019	-73.291	1	36.1	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	CT00-0047-A	03-AUG-2000	41.102	-72.934	1	22.6	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	CT00-0049-A	29-AUG-2000	41.234	-72.265	1	36.9	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	CT00-0053-A	04-AUG-2000	41.328	-71.869	1	1.2	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	CT00-0055-A	19-SEP-2000	41.097	-73.166	1	11.3	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	CT00-0057-A	18-SEP-2000	41.126	-72.965	1	18.3	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	CT00-0059-A	18-SEP-2000	41.164	-72.924	1	17.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	CT00-0061-A	19-SEP-2000	41.203	-72.998	1	9.1	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	CT00-0063-A	19-SEP-2000	41.225	-72.965	1	8.2	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	CT00-0065-A	25-SEP-2000	41.235	-72.815	1	10.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	CT00-0067-A	25-SEP-2000	41.248	-72.577	1	11.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	CT00-0069-A	07-SEP-2000	41.243	-72.335	1	9.1	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0002-A	26-SEP-2001	41.176	-73.123	1	1.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0004-B	26-SEP-2001	41.248	-72.927	1	3.2	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0006-A	21-SEP-2001	41.309	-73.077	1	1.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0008-A	26-SEP-2001	41.28	-72.909	1	1.6	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0010-A	19-SEP-2001	41.28	-72.318	1	3.2	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0012-A	27-SEP-2001	41.325	-71.97	1	1.6	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0014-A	19-SEP-2001	41.374	-72.369	1	2.9	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0016-A	28-SEP-2001	41.422	-72.091	1	2.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0018-A	28-SEP-2001	41.472	-72.073	1	1.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0020-A	28-SEP-2001	41.502	-72.085	1	1.5	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0024-A	30-AUG-2001	41.041	-73.418	1	13.9	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0026-A	30-AUG-2001	41.109	-73.253	1	10.5	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0027-A	05-SEP-2001	41.058	-73.234	1	21.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0028-A	01-AUG-2001	41.122	-73.09	1	12.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0030-A	01-AUG-2001	41.082	-73.022	1	25.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0031-A	06-SEP-2001	41.164	-73.014	1	12.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0032-A	29-AUG-2001	41.159	-72.849	1	19.1	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0033-A	06-SEP-2001	41.14	-72.948	1	18.4	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0034-A	06-SEP-2001	41.232	-72.829	1	9.3	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0036-A	10-SEP-2001	41.271	-72.275	1	7.1	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0038-A	07-AUG-2001	41.071	-73.336	1	8.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0040-A	30-AUG-2001	40.994	-73.411	1	41.8	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0042-A	01-AUG-2001	41.08	-73.165	1	19.4	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0043-A	30-AUG-2001	40.984	-73.502	1	32.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0044-A	06-AUG-2001	41.178	-72.96	1	14.5	m	
National Coastal Assessment-Northeast/University of Rhode Island	2001	CT01-0046-A	18-JUL-2001	41.312	-71.991	1	3.3	m	
National Coastal Assessment-Northeast/University of Rhode Island	2001	CT01-0048-A	18-JUL-2001	41.339	-71.976	1	1.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0050-A	12-SEP-2001	41.247	-72.331	1	8.2	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0052-A	12-SEP-2001	41.236	-72.404	1	11.6	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0054-A	14-SEP-2001	41.244	-72.574	1	9.8	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0056-A	14-SEP-2001	41.207	-72.719	1	12.2	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0058-A	18-SEP-2001	41.077	-72.759	1	29.9	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0060-A	17-SEP-2001	41.1	-72.663	1	26.8	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0062-A	24-SEP-2001	41.007	-73.505	1	21.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0064-A	21-SEP-2001	41.076	-73.078	1	19.8	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0066-A	21-SEP-2001	41.062	-73.265	1	19.5	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0068-A	24-SEP-2001	40.957	-73.41	1	13.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0070-A	26-SEP-2001	40.942	-73.637	1	17.6	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	CT01-0072-A	27-SEP-2001	41.232	-73.012	1	9.1	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	CT02-0200-A	18-SEP-2002	41.146	-73.217	1	3.3	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	CT02-0202-A	28-AUG-2002	41.225	-73.112	1	1.8	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	CT02-0203-A	18-SEP-2002	41.274	-72.927	1	2.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	CT02-0205-A	28-AUG-2002	41.31	-73.079	1	2.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	CT02-0206-A	28-AUG-2002	41.299	-73.066	1	7.8	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	CT02-0207-A	18-SEP-2002	41.286	-72.909	1	8.1	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	CT02-0208-A	24-SEP-2002	41.332	-72.344	1	1.8	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	CT02-0210-A	25-SEP-2002	41.319	-72.086	1	7.1	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	CT02-0212-A	24-SEP-2002	41.403	-72.41	1	3.9	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	CT02-0213-A	24-SEP-2002	41.383	-72.355	1	3.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	CT02-0215-A	25-SEP-2002	41.413	-72.093	1	4.5	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	CT02-0217-A	25-SEP-2002	41.452	-72.081	1	1.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	CT02-0219-A	25-SEP-2002	41.504	-72.086	1	5.2	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	CT02-0220-A	01-OCT-2002	41.002	-73.481	1	23.5	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	CT02-0221-A	24-SEP-2002	41.029	-73.317	1	21.6	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	CT02-0222-A	24-SEP-2002	41.039	-73.364	1	16.2	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	CT02-0223-A	24-SEP-2002	41.088	-73.31	1	12.1	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	CT02-0224-A	24-SEP-2002	41.085	-73.178	1	16.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	CT02-0225-A	25-SEP-2002	41.101	-73.32	1	12.8	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	CT02-0226-A	25-SEP-2002	41.176	-73.016	1	9.1	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	CT02-0227-A	20-SEP-2002	41.193	-72.695	1	20.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	CT02-0228-A	23-SEP-2002	41.232	-72.967	1	8.2	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	CT02-0229-A	17-SEP-2002	41.232	-72.396	1	8.2	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	CT02-0230-A	17-SEP-2002	41.233	-72.403	1	9.8	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	CT02-0231-A	17-SEP-2002	41.245	-72.255	1	33.2	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	CT02-0232-A	17-SEP-2002	41.236	-72.285	1	32.6	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	CT02-0233-A	16-SEP-2002	41.289	-72.199	1	7.9	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	CT02-0234-A	16-SEP-2002	41.318	-72.083	1	8.2	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2003	CT03-0021-A	20-AUG-2003	40.963	-73.623	1	14.1	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2003	CT03-0034-A	27-AUG-2003	41.232	-72.829	1	10.1	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2003	CT03-0035-A	27-AUG-2003	41.209	-72.908	1	11.1	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2003	CT03-0039-A	27-AUG-2003	41.242	-72.665	1	10.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2003	CT03-0241-A	22-SEP-2003	41.132	-72.841	1	25.3	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2003	CT03-0242-A	15-SEP-2003	41.15	-72.695	1	28.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2003	CT03-0243-A	26-SEP-2003	41.181	-73.055	1	9.1	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2003	CT03-0244-A	17-SEP-2003	41.194	-72.78	1	14.6	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2003	CT03-0245-A	17-SEP-2003	41.247	-72.582	1	7.9	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2004	CT04-0023-A	03-SEP-2004	40.979	-73.56	1	21.9	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2004	CT04-0027-A	20-AUG-2004	41.058	-73.234	1	20.8	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2004	CT04-0029-A	07-SEP-2004	41.12	-73.162	1	9.5	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2004	CT04-0030-A	07-SEP-2004	41.082	-73.022	1	25.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2004	CT04-0032-A	19-AUG-2004	41.159	-72.849	1	20.8	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2004	CT04-0040-A	03-SEP-2004	40.994	-73.411	1			
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2004	CT04-0044-A	07-SEP-2004	41.178	-72.96	1	13.4	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2004	CT04-0049-A	19-JUL-2004	41.234	-72.265	1	36.2	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2004	CT04-0223-A	27-SEP-2004	41.088	-73.312	1	11.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2004	CT04-0309-A	24-SEP-2004	41.27	-72.926	1	2.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2004	CT04-0312-A	17-SEP-2004	41.332	-72.18	1	1.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2004	CT04-0313-A	22-SEP-2004	41.324	-71.97	1	2.1	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2004	CT04-0316-A	20-SEP-2004	41.428	-72.1	1	1.9	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2004	CT04-0317-A	22-SEP-2004	41.348	-71.97	1			
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2004	CT04-0401-A	27-SEP-2004	41.057	-73.221	1	22.6	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2004	CT04-0402-A	22-SEP-2004	41.117	-72.965	1	22.6	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2004	CT04-0404-A	20-SEP-2004	41.185	-72.92	1	14.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2004	CT04-0405-A	20-SEP-2004	41.238	-72.726	1	7.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2005	CT05-0001-A	22-SEP-2005	41.241	-72.932	1	3.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2005	CT05-0003-A	19-SEP-2005	41.018	-73.144	1	40.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2005	CT05-0004-A	21-JUL-2005	41.058	-73.234	1	22.1	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2005	CT05-0008-A	22-SEP-2005	41.242	-72.665	1	11.6	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2005	CT05-0011-A	23-SEP-2005	41.551	-72.557	1	2.8	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2005	CT05-0012-A	19-SEP-2005	40.994	-73.411	1	43.9	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2005	CT05-0013-A	15-SEP-2005	40.961	-73.476	1	14.2	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2005	CT05-0015-A	19-SEP-2005	41.009	-73.513	1	14.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2005	CT05-0017-A	26-SEP-2005	41.28	-72.364	1	5.5	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2005	CT05-0018-A	07-JUL-2005	41.055	-73.08	1	25.3	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2005	CT05-0019-A	15-SEP-2005	40.956	-73.58	1	20.4	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2005	CT05-0021-A	15-SEP-2005	40.873	-73.734	1	32.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2005	CT05-0023-A	07-JUL-2005	41.138	-72.655	1	27.6	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2005	CT05-0024-A	19-SEP-2005	41.019	-73.291	1	37.8	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2005	CT05-0025-A	22-SEP-2005	41.178	-72.96	1	15.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2005	CT05-0051-A	28-SEP-2005	41.016	-73.455	1		m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2005	CT05-0052-A	13-SEP-2005	41.046	-72.642	1		m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2005	CT05-0053-A	30-SEP-2005	41.075	-73.26	1		m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2005	CT05-0054-A	19-SEP-2005	41.095	-72.869	1		m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2005	CT05-0055-A	19-SEP-2005	41.124	-72.927	1		m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2005	CT05-0056-A	14-SEP-2005	41.148	-72.484	1		m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2005	CT05-0057-A	15-SEP-2005	41.17	-72.533	1		m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2005	CT05-0058-A	09-SEP-2005	41.222	-72.248	1		m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2005	CT05-0059-A	08-SEP-2005	41.243	-72.335	1		m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2005	CT05-0060-A	09-SEP-2005	41.291	-72.172	1		m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2005	CT05-0061-A	28-SEP-2005	40.933	-73.543	1		m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0002-A	13-SEP-2006	41.078	-72.833	1	29.6	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0003-A	03-AUG-2006	41.018	-73.144	1	39.3	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0005-A	01-AUG-2006	41.237	-72.053	1	72.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0006-A	14-AUG-2006	41.246	-72.468	1	12.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0007-A	07-AUG-2006	41.004	-72.651	1	20.1	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0009-A	03-OCT-2006	41.12	-73.162	1	11.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0010-A	03-OCT-2006	41.122	-73.09	1	13.4	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0014-A	01-AUG-2006	41.026	-72.913	1	40.1	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0014-A	16-AUG-2006	41.026	-72.913	1	38.8	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0016-A	16-AUG-2006	40.981	-72.918	1	9.8	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0020-A	13-SEP-2006	41.14	-72.948	1	19.3	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0022-A	21-SEP-2006	41.109	-73.253	1	10.3	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0026-A	14-SEP-2006	41.343	-72.365	1	1.9	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0027-A	16-AUG-2006	41.004	-72.768	1	24.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0028-A	02-AUG-2006	40.935	-73.6	1	14.1	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0029-A	03-AUG-2006	41.08	-73.165	1	19.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0030-A	27-JUL-2006	40.984	-73.502	1	31.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0031-A	01-AUG-2006	41.102	-72.934	1	24.4	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0031-A	21-AUG-2006	41.102	-72.934	1	24.4	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0032-A	14-SEP-2006	41.442	-72.457	1	3.2	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0033-A	07-AUG-2006	40.994	-73.042	1	23.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0033-A	18-AUG-2006	40.994	-73.042	1	21.4	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0034-A	21-SEP-2006	41.071	-73.336	1	10.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0035-A	03-AUG-2006	41.082	-73.022	1	26.8	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0036-A	12-SEP-2006	41.196	-72.775	1	15.2	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0037-A	27-JUL-2006	40.963	-73.623	1	16.1	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0038-A	18-SEP-2006	41.384	-72.095	1	2.3	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0039-A	28-SEP-2006	40.952	-73.332	1	16.9	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0040-A	13-SEP-2006	41.209	-72.908	1	11.3	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0041-A	19-SEP-2006	41.273	-72.906	1	2.2	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0042-A	12-SEP-2006	41.232	-72.829	1	11.2	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0043-A	28-SEP-2006	40.95	-73.425	1	12.2	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0045-A	07-AUG-2006	41.098	-72.45	1	20.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0047-A	04-AUG-2006	41.164	-73.014	1	14.9	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0048-A	28-SEP-2006	41.041	-73.418	1	12.2	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0049-A	14-AUG-2006	41.271	-72.275	1	6.6	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0050-A	27-JUL-2006	40.979	-73.56	1	24.2	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0075-A	04-OCT-2006	41.016	-73.455	1		m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0076-A	10-OCT-2006	41.018	-73.226	1		m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0077-A	03-OCT-2006	41.04	-72.993	1		m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0078-A	03-OCT-2006	41.094	-73.128	1		m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0079-A	12-OCT-2006	41.057	-73.305	1		m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0080-A	11-SEP-2006	41.205	-72.715	1		m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0081-A	11-SEP-2006	41.247	-72.607	1		m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0082-A	07-SEP-2006	41.061	-72.631	1		m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0083-A	07-SEP-2006	41.161	-72.433	1		m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2006	CT06-0084-A	06-SEP-2006	41.229	-72.402	1		m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DB05-0001-A	04-AUG-2005	39.123	-75.347	1	4.2	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DB05-0003-A	08-AUG-2005	39.537	-75.767	1	12.9	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DB05-0004-A	30-JUL-2005	39.083	-75.183	1	15.0	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DB05-0005-A	05-AUG-2005	38.797	-75.114	1	3.3	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DB05-0006-A	30-JUL-2005	39.093	-75.064	1	4.7	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DB05-0007-A	18-AUG-2005	38.899	-75.179	1	3.2	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DB05-0008-A	26-JUL-2005	38.899	-75.004	1	8.9	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DB05-0009-A	11-AUG-2005	39.216	-75.196	1	3.5	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DB05-0010-B	28-JUL-2005	39.181	-75.107	1	1.3	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DB05-0011-A	01-AUG-2005	39.845	-75.338	1	10.7	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DB05-0012-A	09-AUG-2005	38.931	-75.248	1	3.3	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DB05-0013-A	29-JUL-2005	38.97	-75.202	1	17.0	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DB05-0014-A	11-AUG-2005	39.164	-75.17	1	4.0	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DB05-0015-B	27-JUL-2005	39.107	-75.005	1	3.8	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DB05-0016-A	01-AUG-2005	39.983	-75.067	1	11.0	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DB05-0018-A	28-JUL-2005	39.225	-75.03	1	6.3	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DB05-0019-A	31-JUL-2005	39.653	-75.546	1	10.6	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DB05-0020-A	27-JUL-2005	38.97	-74.967	1	1.2	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DB05-0021-A	08-AUG-2005	39.542	-75.691	1	12.6	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DB05-0022-A	31-JUL-2005	39.374	-75.468	1	7.1	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DB05-0023-A	04-AUG-2005	39.252	-75.364	1	6.0	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DB05-0024-A	29-JUL-2005	39.068	-75.221	1	14.0	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DB06-0002-A	06-SEP-2006	39.389	-75.319	1	1.6	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DB06-0017-A	07-SEP-2006	39.646	-75.461	1	1.0	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DB06-0025-A	07-SEP-2006	39.611	-75.463	1	1.9	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DB06-0026-A	14-AUG-2006	39.704	-75.615	1	0.9	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DB06-0027-A	24-AUG-2006	39.218	-75.044	1	1.7	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DB06-0028-A	03-AUG-2006	39.083	-75.183	1	13.0	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DB06-0028-A	04-AUG-2006	39.083	-75.183	2	12.0	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DB06-0029-A	05-AUG-2006	39.155	-75.064	1	2.1	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DB06-0030-B	07-SEP-2006	39.593	-75.469	1	1.3	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DB06-0031-A	10-AUG-2006	39.269	-75.238	1	3.2	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DB06-0032-A	06-SEP-2006	39.416	-75.417	1	1.9	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DB06-0033-A	08-AUG-2006	39.053	-75.327	1	3.5	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DB06-0034-A	23-AUG-2006	39.574	-75.545	1	8.2	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DB06-0035-C	24-AUG-2006	39.196	-74.897	1	1.9	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DB06-0036-A	25-AUG-2006	39.983	-75.067	1	5.8	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DB06-0037-A	01-AUG-2006	39.073	-75.021	1	2.9	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DB06-0038-A	16-AUG-2006	39.408	-75.6	1	3.1	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DB06-0039-A	10-AUG-2006	39.287	-75.236	1	4.0	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DB06-0040-C	07-SEP-2006	39.614	-75.444	1	1.8	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DB06-0041-A	04-AUG-2006	39.033	-75.255	1	12.0	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DB06-0042-A	23-AUG-2006	39.653	-75.546	1	11.3	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DB06-0043-A	14-AUG-2006	39.501	-75.533	1	0.8	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DB06-0044-A	03-AUG-2006	39.374	-75.468	1	13.0	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DB06-0045-A	24-AUG-2006	39.3	-74.984	1	1.9	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DB06-0046-A	02-AUG-2006	38.814	-75.097	1	21.0	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DB06-0047-A	05-AUG-2006	39.069	-75.155	1	5.4	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DB06-0048-A	09-AUG-2006	38.86	-75.205	1	3.2	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DB06-0049-B	08-SEP-2006	39.835	-75.337	1	0.8	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DB06-0050-A	08-AUG-2006	39.158	-75.392	1	2.8	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2000	DE00-0001-A	17-OCT-2000	38.452	-75.078	1	1.7	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2000	DE00-0003-A	17-OCT-2000	38.485	-75.103	1	0.7	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2000	DE00-0005-A	11-OCT-2000	38.546	-75.199	1	0.7	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2000	DE00-0007-A	19-OCT-2000	38.573	-75.673	1	0.7	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2000	DE00-0009-A	10-OCT-2000	38.564	-75.204	1	1.1	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2000	DE00-0011-B	16-OCT-2000	38.551	-75.101	1	1.6	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2000	DE00-0013-A	20-OCT-2000	38.589	-75.662	1	0.9	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2000	DE00-0015-A	12-OCT-2000	38.594	-75.284	1	1.0	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2000	DE00-0017-A	12-OCT-2000	38.591	-75.177	1	1.8	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2000	DE00-0019-A	16-OCT-2000	38.596	-75.079	1	1.2	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2000	DE00-0021-A	20-OCT-2000	38.615	-75.639	1	1.5	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2000	DE00-0023-A	20-OCT-2000	38.643	-75.571	1	1.3	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2000	DE00-0025-A	18-OCT-2000	38.635	-75.121	1	1.9	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2000	DE00-0027-B	20-OCT-2000	38.644	-75.579	1	1.4	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2000	DE00-0029-A	18-OCT-2000	38.67	-75.127	1	1.3	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2000	DE00-0031-A	18-OCT-2000	38.669	-75.073	1	0.6	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2000	DE00-0033-A	18-OCT-2000	38.685	-75.101	1	1.9	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2000	DE00-0035-B	19-OCT-2000	38.712	-75.179	1	0.5	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	DE00-0037-A	28-SEP-2000	39.225	-75.401	1	3.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	DE00-0039-A	09-OCT-2000	39.063	-75.381	1	1.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	DE00-0041-A	10-OCT-2000	38.995	-75.293	1	5.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	DE00-0043-A	02-OCT-2000	38.864	-75.223	1	3.5	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	DE00-0045-A	02-OCT-2000	38.8	-75.134	1	6.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	DE00-0047-A	11-OCT-2000	39.767	-75.474	1	15.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	DE00-0049-A	11-OCT-2000	39.653	-75.546	1	13.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	DE00-0051-A	05-OCT-2000	39.511	-75.553	1	14.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	DE00-0053-A	04-OCT-2000	39.374	-75.468	1	15.5	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	DE00-0055-A	10-OCT-2000	39.204	-75.359	1	3.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	DE00-0057-A	03-OCT-2000	38.917	-75.1	1	13.4	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	DE00-0059-A	27-SEP-2000	38.797	-75.246	1	3.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	DE00-0061-A	28-SEP-2000	39.244	-75.451	1	4.1	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	DE00-0065-B	29-SEP-2000	39.392	-75.54	1	2.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	DE00-0067-A	06-OCT-2000	39.534	-75.774	1	9.1	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	DE00-0069-B	22-SEP-2000	39.736	-75.535	1	4.5	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2001	DE01-0002-A	18-SEP-2001	38.474	-75.072	1	1.6	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2001	DE01-0004-A	18-SEP-2001	38.485	-75.069	1	0.9	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2001	DE01-0006-A	17-SEP-2001	38.559	-75.698	1	1.9	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2001	DE01-0008-A	17-SEP-2001	38.564	-75.628	1	1.5	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2001	DE01-0010-A	19-SEP-2001	38.568	-75.185	1	1.8	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2001	DE01-0012-A	20-SEP-2001	38.565	-75.094	1	0.6	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2001	DE01-0014-A	01-OCT-2001	38.604	-75.654	1	1.8	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2001	DE01-0016-A	19-SEP-2001	38.591	-75.243	1	1.9	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2001	DE01-0018-A	19-SEP-2001	38.586	-75.149	1	0.5	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2001	DE01-0020-A	20-SEP-2001	38.584	-75.067	1	1.3	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2001	DE01-0022-A	01-OCT-2001	38.634	-75.616	1	1.8	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2001	DE01-0024-A	19-SEP-2001	38.615	-75.161	1	0.9	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2001	DE01-0026-A	20-SEP-2001	38.631	-75.082	1	1.1	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2001	DE01-0028-A	02-OCT-2001	38.664	-75.177	1	1.6	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2001	DE01-0030-A	20-SEP-2001	38.653	-75.101	1	1.9	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2001	DE01-0032-A	03-OCT-2001	38.71	-75.174	1	0.4	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2001	DE01-0034-A	03-OCT-2001	38.687	-75.081	1	1.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	DE01-0036-A	01-AUG-2001	39.244	-75.402	1	2.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	DE01-0038-A	01-AUG-2001	39.231	-75.395	1	1.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	DE01-0040-A	04-OCT-2001	39.08	-75.277	1	8.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	DE01-0042-A	05-OCT-2001	38.932	-75.187	1	9.4	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	DE01-0044-A	05-OCT-2001	38.876	-75.132	1	20.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	DE01-0046-A	10-OCT-2001	39.798	-75.426	1	14.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	DE01-0048-A	10-OCT-2001	39.718	-75.506	1	14.1	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	DE01-0050-A	07-OCT-2001	39.589	-75.563	1	14.5	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	DE01-0052-A	07-OCT-2001	39.453	-75.56	1	12.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	DE01-0054-A	06-OCT-2001	39.3	-75.382	1	14.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	DE01-0056-A	04-OCT-2001	39.167	-75.283	1	12.1	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	DE01-0058-A	31-JUL-2001	38.953	-75.322	1	3.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	DE01-0060-A	31-JUL-2001	39.048	-75.394	1	3.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	DE01-0062-A	02-AUG-2001	39.07	-75.415	1	3.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	DE01-0064-A	01-AUG-2001	39.244	-75.566	1	2.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	DE01-0066-A	30-JUL-2001	39.345	-75.499	1	0.4	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	DE01-0068-A	30-JUL-2001	39.461	-75.638	1	3.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	DE01-0070-A	12-OCT-2001	39.544	-75.673	1	12.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	DE01-0072-A	11-OCT-2001	39.72	-75.519	1	11.5	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	DE01-0074-A	21-AUG-2001	39.736	-75.557	2	4.5	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2001	DE01-0075-A	03-OCT-2001	38.698	-75.096	1	0.7	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2001	DE01-0076-A	02-OCT-2001	38.657	-75.181	1	1.8	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2001	DE01-0077-A	02-OCT-2001	38.636	-75.166	1	0.7	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2001	DE01-0078-A	28-SEP-2001	38.505	-75.094	1	0.8	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2002	DE02-0009-A	02-OCT-2002	38.564	-75.204	1	0.5	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2002	DE02-0021-A	19-SEP-2002	38.615	-75.639	1	1.5	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2002	DE02-0033-A	11-SEP-2002	38.685	-75.102	1	1.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	DE02-0047-A	07-AUG-2002	39.767	-75.474	1	14.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	DE02-0049-A	07-AUG-2002	39.653	-75.546	1	14.5	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	DE02-0051-A	01-AUG-2002	39.511	-75.553	1	14.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	DE02-0053-A	01-AUG-2002	39.374	-75.468	1	13.8	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	DE02-0055-A	31-JUL-2002	39.204	-75.359	1	3.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	DE02-0055-A	01-AUG-2002	39.204	-75.359	2	3.1	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	DE02-0057-A	29-JUL-2002	38.917	-75.1	1	14.8	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2002	DE02-0200-B	26-SEP-2002	38.454	-75.087	1	0.9	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2002	DE02-0202-A	26-SEP-2002	38.482	-75.116	1	1.1	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2002	DE02-0204-C	02-OCT-2002	38.563	-75.192	1	0.4	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2002	DE02-0205-A	12-SEP-2002	38.558	-75.695	1	0.6	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2002	DE02-0207-A	12-SEP-2002	38.565	-75.632	1	1.0	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2002	DE02-0209-A	03-OCT-2002	38.551	-75.101	1	1.0	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2002	DE02-0211-A	12-SEP-2002	38.585	-75.669	1	0.6	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2002	DE02-0213-A	01-OCT-2002	38.593	-75.283	1	0.9	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2002	DE02-0215-A	01-OCT-2002	38.589	-75.197	1	1.6	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2002	DE02-0217-A	03-OCT-2002	38.592	-75.107	1	1.7	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2002	DE02-0219-A	19-SEP-2002	38.623	-75.625	1	1.7	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2002	DE02-0222-A	08-OCT-2002	38.64	-75.129	1	1.6	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2002	DE02-0226-A	08-OCT-2002	38.653	-75.151	1	0.9	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2002	DE02-0228-A	09-OCT-2002	38.661	-75.073	1	0.5	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2002	DE02-0231-A	09-OCT-2002	38.712	-75.181	1	0.6	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2002	DE02-0233-A	10-OCT-2002	38.759	-75.111	1	2.0	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2002	DE02-0235-A	11-SEP-2002	38.78	-75.15	1	3.5	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	DE02-0237-A	22-AUG-2002	39.225	-75.401	1	2.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	DE02-0239-A	31-JUL-2002	39.1	-75.314	1	2.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	DE02-0241-A	23-AUG-2002	39.016	-75.311	1	4.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	DE02-0243-A	29-JUL-2002	38.911	-75.214	1	7.8	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	DE02-0245-A	21-AUG-2002	38.801	-75.133	1	5.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	DE02-0246-A	21-AUG-2002	38.804	-75.19	1	3.4	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	DE02-0251-A	22-AUG-2002	39.265	-75.445	1	1.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	DE02-0252-B	20-AUG-2002	39.354	-75.543	1	2.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	DE02-0255-A	17-SEP-2002	39.5	-75.528	1	2.4	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	DE02-0256-A	07-AUG-2002	39.542	-75.727	1	12.8	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	DE02-0259-A	16-SEP-2002	39.736	-75.534	1	0.4	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2003	DE03-0004-A	17-JUL-2003	38.485	-75.069	1	0.8	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2003	DE03-0018-A	16-JUL-2003	38.586	-75.149	1	1.0	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2003	DE03-0034-A	06-AUG-2003	38.687	-75.081	1	1.8	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	DE03-0046-A	06-AUG-2003	39.798	-75.426	1	15.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	DE03-0048-A	06-AUG-2003	39.718	-75.506	1	13.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	DE03-0050-A	31-JUL-2003	39.589	-75.563	1	14.8	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	DE03-0052-A	30-JUL-2003	39.453	-75.56	1	14.4	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	DE03-0052-A	31-JUL-2003	39.453	-75.56	2	11.4	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	DE03-0054-A	30-JUL-2003	39.3	-75.382	1	15.5	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	DE03-0056-A	29-JUL-2003	39.167	-75.283	1	10.8	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2003	DE03-0201-A	17-JUL-2003	38.478	-75.059	1	1.4	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2003	DE03-0205-A	15-JUL-2003	38.558	-75.695	1	1.1	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2003	DE03-0207-A	15-JUL-2003	38.565	-75.632	1	1.4	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2003	DE03-0208-A	16-JUL-2003	38.572	-75.18	1	1.5	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2003	DE03-0210-B	04-AUG-2003	38.555	-75.095	1	0.6	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2003	DE03-0212-A	15-JUL-2003	38.605	-75.653	1	1.6	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2003	DE03-0214-A	16-JUL-2003	38.588	-75.261	1	0.5	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2003	DE03-0218-C	04-AUG-2003	38.586	-75.065	1	0.8	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2003	DE03-0219-A	15-JUL-2003	38.623	-75.625	1	1.9	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2003	DE03-0221-A	16-JUL-2003	38.615	-75.162	1	0.6	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2003	DE03-0223-A	04-AUG-2003	38.623	-75.089	1	1.1	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2003	DE03-0225-A	06-AUG-2003	38.663	-75.175	1	1.2	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2003	DE03-0227-A	05-AUG-2003	38.673	-75.111	1	1.8	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2003	DE03-0229-A	05-AUG-2003	38.698	-75.157	1	0.5	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2003	DE03-0232-A	07-AUG-2003	38.715	-75.093	1	0.9	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2003	DE03-0234-A	07-AUG-2003	38.75	-75.1	1	0.4	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	DE03-0236-A	25-SEP-2003	39.244	-75.403	1	4.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	DE03-0238-A	25-SEP-2003	39.231	-75.395	1	3.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	DE03-0240-A	29-JUL-2003	39.08	-75.276	1	8.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	DE03-0242-A	28-JUL-2003	38.932	-75.186	1	8.5	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	DE03-0244-A	28-JUL-2003	38.877	-75.131	1	19.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	DE03-0247-A	23-SEP-2003	38.946	-75.339	1	2.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	DE03-0248-A	24-SEP-2003	39.066	-75.403	1	4.8	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	DE03-0249-A	24-SEP-2003	39.07	-75.415	1	3.1	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	DE03-0250-A	25-SEP-2003	39.249	-75.479	1	2.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	DE03-0253-A	26-SEP-2003	39.302	-75.476	1	1.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	DE03-0254-B	02-OCT-2003	39.456	-75.649	1	3.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	DE03-0257-A	31-JUL-2003	39.559	-75.574	1	2.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	DE03-0258-A	03-OCT-2003	39.736	-75.557	1	7.9	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2004	DE04-0004-A	08-JUL-2004	38.485	-75.069	1	1.3	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2004	DE04-0009-A	12-JUL-2004	38.564	-75.204	1	0.3	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2004	DE04-0021-A	07-JUL-2004	38.615	-75.639	1	0.6	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2004	DE04-0033-A	09-JUL-2004	38.685	-75.102	1	1.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	DE04-0047-A	11-AUG-2004	39.767	-75.474	1	9.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	DE04-0051-A	05-AUG-2004	39.511	-75.553	1	13.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	DE04-0055-A	04-AUG-2004	39.204	-75.359	1	3.1	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	DE04-0057-A	02-AUG-2004	38.917	-75.1	1	13.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	DE04-0239-A	15-JUL-2004	39.1	-75.314	1	3.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	DE04-0246-A	12-JUL-2004	38.804	-75.19	1	3.1	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	DE04-0254-A	14-JUL-2004	39.456	-75.649	1	1.3	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2004	DE04-0400-A	08-JUL-2004	38.46	-75.084	1	0.5	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2004	DE04-0402-A	08-JUL-2004	38.483	-75.118	1	0.7	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2004	DE04-0403-A	12-JUL-2004	38.548	-75.198	1	0.3	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2004	DE04-0405-A	14-JUL-2004	38.57	-75.64	1	0.6	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2004	DE04-0408-A	13-JUL-2004	38.551	-75.102	1	0.4	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2004	DE04-0410-A	14-JUL-2004	38.589	-75.665	1	0.4	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2004	DE04-0412-B	12-JUL-2004	38.586	-75.275	1	0.8	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2004	DE04-0414-A	12-JUL-2004	38.588	-75.214	1	0.5	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2004	DE04-0415-A	13-JUL-2004	38.601	-75.097	1	1.5	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2004	DE04-0418-A	07-JUL-2004	38.644	-75.571	1	1.0	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2004	DE04-0420-A	09-JUL-2004	38.644	-75.116	1	1.6	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2004	DE04-0422-A	07-JUL-2004	38.645	-75.59	1	1.5	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2004	DE04-0425-A	09-JUL-2004	38.652	-75.074	1	0.3	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2004	DE04-0428-A	09-JUL-2004	38.712	-75.18	1	0.3	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2004	DE04-0430-A	15-JUL-2004	38.774	-75.134	1	1.8	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2004	DE04-0432-A	15-JUL-2004	38.779	-75.143	1	0.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	DE04-0434-A	13-JUL-2004	39.151	-75.405	1	1.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	DE04-0437-A	13-JUL-2004	39.013	-75.311	1	3.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	DE04-0438-A	02-AUG-2004	38.931	-75.193	1	9.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	DE04-0440-A	12-JUL-2004	38.794	-75.136	1	3.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	DE04-0444-A	15-JUL-2004	39.251	-75.547	1	0.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	DE04-0450-B	09-AUG-2004	39.554	-75.645	1	14.1	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	DE04-0455-A	05-AUG-2004	39.622	-75.6	1	7.2	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DI05-0001-A	22-JUL-2005	38.658	-75.102	1	2.0	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DI05-0002-A	18-JUL-2005	38.691	-75.14	1	0.8	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DI05-0003-B	19-JUL-2005	38.586	-75.156	1	0.9	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DI05-0004-A	22-JUL-2005	38.65	-75.099	1	1.9	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DI05-0005-A	21-JUL-2005	38.621	-75.068	1	0.5	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DI05-0006-A	02-AUG-2005	38.687	-75.081	1	1.6	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DI05-0007-A	21-JUL-2005	38.6	-75.091	1	4.1	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DI05-0008-A	18-JUL-2005	38.463	-75.063	1	1.0	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DI05-0009-A	22-JUL-2005	38.658	-75.094	1	2.0	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DI05-0010-A	18-JUL-2005	38.681	-75.099	1	1.9	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DI05-0011-A	18-JUL-2005	38.588	-75.183	1	1.5	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DI05-0012-A	02-AUG-2005	38.667	-75.115	1	1.7	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DI05-0013-A	18-JUL-2005	38.607	-75.127	1	2.0	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DI05-0014-A	18-JUL-2005	38.493	-75.058	1	0.7	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DI05-0015-A	21-JUL-2005	38.625	-75.078	1	0.3	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DI05-0016-A	20-JUL-2005	38.506	-75.071	1	0.6	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DI05-0017-A	18-JUL-2005	38.592	-75.282	1	0.7	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DI05-0018-A	19-JUL-2005	38.613	-75.103	1	0.9	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DI05-0019-A	19-JUL-2005	38.607	-75.137	1	2.0	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DI05-0020-A	20-JUL-2005	38.48	-75.079	1	1.4	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DI05-0021-A	22-SEP-2005	38.642	-75.136	1	0.5	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DI05-0022-A	03-AUG-2005	38.64	-75.128	1	1.7	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DI05-0023-A	18-JUL-2005	38.576	-75.183	1	1.3	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DI05-0024-A	18-JUL-2005	38.667	-75.098	1	1.9	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2005	DI05-0025-A	18-JUL-2005	38.593	-75.208	1	1.9	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DI06-0026-A	26-SEP-2006	38.586	-75.669	1	0.5	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DI06-0027-A	11-JUL-2006	38.608	-75.079	1	4.2	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DI06-0028-A	07-JUL-2006	38.602	-75.114	1	1.8	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DI06-0029-A	05-JUL-2006	38.457	-75.086	1	1.1	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DI06-0030-A	06-JUL-2006	38.607	-75.151	1	1.2	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DI06-0031-A	17-JUL-2006	38.693	-75.107	1	0.9	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DI06-0032-A	06-JUL-2006	38.579	-75.167	1	1.4	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DI06-0033-A	18-JUL-2006	38.657	-75.115	1	2.3	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DI06-0034-A	06-JUL-2006	38.585	-75.261	1	0.7	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DI06-0035-A	17-JUL-2006	38.69	-75.079	1	0.9	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DI06-0036-A	11-JUL-2006	38.582	-75.096	1	2.4	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DI06-0037-A	05-JUL-2006	38.479	-75.073	1	1.4	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DI06-0038-A	07-JUL-2006	38.595	-75.123	1	1.3	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DI06-0039-A	12-JUL-2006	38.645	-75.106	1	1.5	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DI06-0040-A	12-JUL-2006	38.656	-75.173	1	0.6	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DI06-0041-A	17-JUL-2006	38.674	-75.092	1	1.9	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DI06-0042-A	12-JUL-2006	38.65	-75.091	1	0.9	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DI06-0043-A	18-JUL-2006	38.684	-75.132	1	1.5	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DI06-0044-A	06-JUL-2006	38.601	-75.168	1	0.3	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DI06-0045-A	18-JUL-2006	38.67	-75.124	1	1.3	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DI06-0046-A	12-JUL-2006	38.634	-75.084	1	1.6	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DI06-0047-A	17-JUL-2006	38.675	-75.081	1	1.9	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DI06-0048-A	07-JUL-2006	38.596	-75.114	1	1.9	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DI06-0049-A	11-JUL-2006	38.568	-75.095	1	1.4	m	
National Coastal Assessment-Northeast/Delaware Dept. of Natural Resources	2006	DI06-0050-A	11-JUL-2006	38.59	-75.085	1	1.3	m	
R-EMAP Region 2 1993-94	1993	JB002	14-SEP-1993	40.636	-73.798	1	2.7	m	
R-EMAP Region 2 1993-94	1993	JB006	16-SEP-1993	40.608	-73.773	1	4.0	m	
R-EMAP Region 2 1993-94	1993	JB008	14-SEP-1993	40.641	-73.816	1	9.4	m	
R-EMAP Region 2 1998	1998	JB008	01-JUL-1998	40.641	-73.816	1			
R-EMAP Region 2 1998	1998	JB008	04-AUG-1998	40.641	-73.816	2	8.8	m	
R-EMAP Region 2 1993-94	1993	JB012	24-SEP-1993	40.648	-73.89	1	3.0	m	
R-EMAP Region 2 1993-94	1993	JB015	15-SEP-1993	40.626	-73.794	1	10.1	m	
R-EMAP Region 2 1993-94	1993	JB018	15-SEP-1993	40.609	-73.786	1	16.2	m	
R-EMAP Region 2 1998	1998	JB018	01-JUL-1998	40.61	-73.786	1			
R-EMAP Region 2 1998	1998	JB018	05-AUG-1998	40.61	-73.786	2	13.4	m	
R-EMAP Region 2 1993-94	1993	JB022	17-SEP-1993	40.604	-73.78	1	2.6	m	
R-EMAP Region 2 1993-94	1993	JB026	16-SEP-1993	40.603	-73.842	1	5.2	m	
R-EMAP Region 2 1998	1998	JB026	01-JUL-1998	40.603	-73.842	1			
R-EMAP Region 2 1998	1998	JB026	07-AUG-1998	40.603	-73.842	2	5.8	m	
R-EMAP Region 2 1993-94	1993	JB031	17-SEP-1993	40.611	-73.872	1	2.7	m	
R-EMAP Region 2 1998	1998	JB031	01-JUL-1998	40.611	-73.872	1			
R-EMAP Region 2 1998	1998	JB031	07-AUG-1998	40.611	-73.872	2			
R-EMAP Region 2 1998	1998	JB031	08-AUG-1998	40.611	-73.872	3	2.7	m	
R-EMAP Region 2 1993-94	1993	JB033	13-SEP-1993	40.616	-73.888	1	12.2	m	
R-EMAP Region 2 1998	1998	JB033	01-JUL-1998	40.616	-73.888	1			
R-EMAP Region 2 1998	1998	JB033	03-AUG-1998	40.616	-73.888	2	12.5	m	
R-EMAP Region 2 1993-94	1993	JB039	08-SEP-1993	40.587	-73.846	1	5.8	m	
R-EMAP Region 2 1998	1998	JB039	01-JUL-1998	40.587	-73.845	1			
R-EMAP Region 2 1998	1998	JB039	01-AUG-1998	40.587	-73.845	2	6.1	m	
R-EMAP Region 2 1993-94	1993	JB041	09-SEP-1993	40.586	-73.86	1	7.9	m	
R-EMAP Region 2 1998	1998	JB041	01-JUL-1998	40.585	-73.861	1			
R-EMAP Region 2 1998	1998	JB041	01-AUG-1998	40.585	-73.861	2	8.2	m	
R-EMAP Region 2 1993-94	1993	JB042	17-SEP-1993	40.583	-73.848	1	7.6	m	
R-EMAP Region 2 1998	1998	JB042	01-JUL-1998	40.583	-73.847	1			
R-EMAP Region 2 1998	1998	JB042	01-AUG-1998	40.583	-73.847	2	6.7	m	
R-EMAP Region 2 1993-94	1993	JB043	09-SEP-1993	40.576	-73.874	1	10.1	m	
R-EMAP Region 2 1998	1998	JB043	01-JUL-1998	40.576	-73.875	1			
R-EMAP Region 2 1998	1998	JB043	17-JUL-1998	40.576	-73.875	2	9.4	m	
R-EMAP Region 2 1993-94	1994	JB101	09-SEP-1994	40.64	-73.814	1	7.6	m	
R-EMAP Region 2 1993-94	1994	JB103	12-SEP-1994	40.629	-73.788	1	6.7	m	
R-EMAP Region 2 1993-94	1994	JB104	12-SEP-1994	40.622	-73.842	1	2.4	m	
R-EMAP Region 2 1993-94	1994	JB106	06-SEP-1994	40.621	-73.89	1	13.4	m	
R-EMAP Region 2 1993-94	1994	JB108	08-SEP-1994	40.617	-73.857	1	2.7	m	
R-EMAP Region 2 1993-94	1994	JB110	09-SEP-1994	40.607	-73.815	1	7.3	m	
R-EMAP Region 2 1993-94	1994	JB111	08-SEP-1994	40.605	-73.791	1	10.4	m	
R-EMAP Region 2 1993-94	1994	JB112	08-SEP-1994	40.603	-73.865	1	4.6	m	
R-EMAP Region 2 1993-94	1994	JB113	06-SEP-1994	40.596	-73.867	1	5.2	m	
R-EMAP Region 2 1993-94	1994	JB114	08-SEP-1994	40.591	-73.851	1	5.2	m	
R-EMAP Region 2 1993-94	1994	JB115	06-SEP-1994	40.634	-73.87	1	2.9	m	
R-EMAP Region 2 1993-94	1994	JB117	14-SEP-1994	40.623	-73.765	1	4.6	m	
R-EMAP Region 2 1993-94	1994	JB119	12-SEP-1994	40.604	-73.875	1	3.1	m	
R-EMAP Region 2 1993-94	1994	JB120	13-SEP-1994	40.596	-73.813	1	3.7	m	
R-EMAP Region 2 1998	1998	JB201	01-JUL-1998	40.572	-73.879	1			
R-EMAP Region 2 1998	1998	JB201	17-JUL-1998	40.572	-73.879	2	11.0	m	
R-EMAP Region 2 1998	1998	JB202	01-JUL-1998	40.612	-73.81	1			
R-EMAP Region 2 1998	1998	JB202	06-AUG-1998	40.612	-73.81	2	4.0	m	
R-EMAP Region 2 1998	1998	JB203	01-JUL-1998	40.633	-73.807	1			
R-EMAP Region 2 1998	1998	JB203	04-AUG-1998	40.633	-73.807	2	11.9	m	
R-EMAP Region 2 1998	1998	JB204	01-JUL-1998	40.608	-73.89	1			
R-EMAP Region 2 1998	1998	JB204	03-AUG-1998	40.608	-73.89	2	9.1	m	
R-EMAP Region 2 1998	1998	JB205	01-JUL-1998	40.589	-73.859	1			
R-EMAP Region 2 1998	1998	JB205	01-AUG-1998	40.589	-73.859	2	2.7	m	
R-EMAP Region 2 1998	1998	JB206	01-JUL-1998	40.595	-73.805	1			
R-EMAP Region 2 1998	1998	JB206	05-AUG-1998	40.595	-73.805	2	5.5	m	
R-EMAP Region 2 1998	1998	JB207	01-JUL-1998	40.629	-73.759	1			
R-EMAP Region 2 1998	1998	JB207	06-AUG-1998	40.629	-73.759	2	7.6	m	
R-EMAP Region 2 1998	1998	JB209	01-JUL-1998	40.605	-73.787	1			
R-EMAP Region 2 1998	1998	JB209	05-AUG-1998	40.605	-73.787	2	9.4	m	
R-EMAP Region 2 1998	1998	JB210	01-JUL-1998	40.628	-73.871	1			
R-EMAP Region 2 1998	1998	JB210	08-AUG-1998	40.628	-73.871	2	2.1	m	
R-EMAP Region 2 1998	1998	JB211	01-JUL-1998	40.612	-73.873	1			
R-EMAP Region 2 1998	1998	JB211	08-AUG-1998	40.612	-73.873	2	2.7	m	
R-EMAP Region 2 1998	1998	JB212	01-JUL-1998	40.588	-73.834	1			
R-EMAP Region 2 1998	1998	JB212	06-AUG-1998	40.588	-73.834	2	2.1	m	
R-EMAP Region 2 1998	1998	JB213	01-JUL-1998	40.619	-73.778	1			
R-EMAP Region 2 1998	1998	JB213	05-AUG-1998	40.619	-73.778	2	10.1	m	
R-EMAP Region 2 1998	1998	JB214	01-JUL-1998	40.643	-73.858	1			
R-EMAP Region 2 1998	1998	JB214	03-AUG-1998	40.643	-73.858	2	6.4	m	
R-EMAP Region 2 1998	1998	JB215	01-JUL-1998	40.626	-73.837	1			
R-EMAP Region 2 1998	1998	JB215	10-AUG-1998	40.626	-73.837	2	3.4	m	
R-EMAP Region 2 1998	1998	JB216	01-JUL-1998	40.633	-73.873	1			
R-EMAP Region 2 1998	1998	JB216	08-AUG-1998	40.633	-73.873	2	11.6	m	
R-EMAP Region 2 1998	1998	JB217	01-JUL-1998	40.585	-73.852	1			
R-EMAP Region 2 1998	1998	JB217	10-AUG-1998	40.585	-73.852	2	9.4	m	
R-EMAP Region 2 1998	1998	JB219	01-JUL-1998	40.575	-73.887	1			
R-EMAP Region 2 1998	1998	JB219	08-AUG-1998	40.575	-73.887	2	10.1	m	
R-EMAP Region 2 1998	1998	JB222	01-JUL-1998	40.603	-73.878	1			
R-EMAP Region 2 1998	1998	JB222	11-AUG-1998	40.603	-73.878	2	8.5	m	
R-EMAP Region 2 1998	1998	JB223	01-JUL-1998	40.593	-73.871	1			
R-EMAP Region 2 1998	1998	JB223	10-AUG-1998	40.593	-73.871	2	11.0	m	
R-EMAP Region 2 2003	2003	JB301	31-JUL-2003	40.629	-73.759	1	9.5	m	
R-EMAP Region 2 2003	2003	JB301	01-AUG-2003	40.629	-73.759	2	9.5	m	
R-EMAP Region 2 2003	2003	JB303	08-AUG-2003	40.619	-73.778	1	10.7	m	
R-EMAP Region 2 2003	2003	JB303	11-AUG-2003	40.619	-73.778	2	10.7	m	
R-EMAP Region 2 2003	2003	JB305	07-AUG-2003	40.575	-73.87	1	4.3	m	
R-EMAP Region 2 2003	2003	JB305	08-AUG-2003	40.575	-73.87	2	4.3	m	
R-EMAP Region 2 2003	2003	JB306	05-AUG-2003	40.572	-73.88	1	5.2	m	
R-EMAP Region 2 2003	2003	JB306	06-AUG-2003	40.572	-73.88	2	5.2	m	
R-EMAP Region 2 2003	2003	JB307	11-AUG-2003	40.64	-73.847	1	6.1	m	
R-EMAP Region 2 2003	2003	JB307	12-AUG-2003	40.64	-73.847	2	6.1	m	
R-EMAP Region 2 2003	2003	JB309	05-AUG-2003	40.643	-73.858	1	12.2	m	
R-EMAP Region 2 2003	2003	JB309	06-AUG-2003	40.643	-73.858	2	12.2	m	
R-EMAP Region 2 2003	2003	JB310	12-AUG-2003	40.639	-73.828	1	1.7	m	
R-EMAP Region 2 2003	2003	JB310	13-AUG-2003	40.639	-73.828	2	1.7	m	
R-EMAP Region 2 2003	2003	JB313	11-AUG-2003	40.61	-73.81	1	10.1	m	
R-EMAP Region 2 2003	2003	JB313	12-AUG-2003	40.61	-73.81	2	10.1	m	
R-EMAP Region 2 2003	2003	JB315	14-AUG-2003	40.605	-73.786	1	2.7	m	
R-EMAP Region 2 2003	2003	JB315	15-AUG-2003	40.605	-73.786	2	2.7	m	
R-EMAP Region 2 2003	2003	JB316	08-AUG-2003	40.625	-73.837	1	11.0	m	
R-EMAP Region 2 2003	2003	JB316	11-AUG-2003	40.625	-73.837	2	11.0	m	
R-EMAP Region 2 2003	2003	JB317	13-AUG-2003	40.621	-73.812	1	7.6	m	
R-EMAP Region 2 2003	2003	JB317	14-AUG-2003	40.621	-73.812	2	7.6	m	
R-EMAP Region 2 2003	2003	JB319	05-AUG-2003	40.633	-73.807	1	10.7	m	
R-EMAP Region 2 2003	2003	JB319	06-AUG-2003	40.633	-73.807	2	10.7	m	
R-EMAP Region 2 2003	2003	JB322	07-AUG-2003	40.627	-73.871	1	6.7	m	
R-EMAP Region 2 2003	2003	JB322	08-AUG-2003	40.627	-73.871	2	6.7	m	
R-EMAP Region 2 2003	2003	JB323	06-AUG-2003	40.633	-73.873	1	11.3	m	
R-EMAP Region 2 2003	2003	JB323	07-AUG-2003	40.633	-73.873	2	11.3	m	
R-EMAP Region 2 2003	2003	JB354	06-AUG-2003	40.602	-73.877	1	11.0	m	
R-EMAP Region 2 2003	2003	JB354	07-AUG-2003	40.602	-73.877	2	11.0	m	
R-EMAP Region 2 2003	2003	JB358	07-AUG-2003	40.608	-73.89	1	7.9	m	
R-EMAP Region 2 2003	2003	JB358	08-AUG-2003	40.608	-73.89	2	7.9	m	
R-EMAP Region 2 2003	2003	JB359	07-AUG-2003	40.612	-73.872	1	3.4	m	
R-EMAP Region 2 2003	2003	JB359	08-AUG-2003	40.612	-73.872	2	3.4	m	
R-EMAP Region 2 2003	2003	JB361	08-AUG-2003	40.584	-73.853	1	3.6	m	
R-EMAP Region 2 2003	2003	JB361	11-AUG-2003	40.584	-73.853	2	3.6	m	
R-EMAP Region 2 2003	2003	JB364	11-AUG-2003	40.593	-73.871	1	5.8	m	
R-EMAP Region 2 2003	2003	JB364	12-AUG-2003	40.593	-73.871	2	5.8	m	
R-EMAP Region 2 2003	2003	JB366	13-AUG-2003	40.589	-73.859	1	4.0	m	
R-EMAP Region 2 2003	2003	JB366	14-AUG-2003	40.589	-73.859	2	4.0	m	
R-EMAP Region 2 2003	2003	JB367	12-AUG-2003	40.588	-73.835	1	7.3	m	
R-EMAP Region 2 2003	2003	JB367	13-AUG-2003	40.588	-73.835	2	7.3	m	
R-EMAP Region 2 2003	2003	JB368	12-AUG-2003	40.592	-73.846	1	5.5	m	
R-EMAP Region 2 2003	2003	JB368	13-AUG-2003	40.592	-73.846	2	5.5	m	
R-EMAP Region 2 2003	2003	JB371	14-AUG-2003	40.595	-73.805	1	7.3	m	
R-EMAP Region 2 2003	2003	JB371	15-AUG-2003	40.595	-73.805	2	7.3	m	
R-EMAP Region 2 2003	2003	JB372	14-AUG-2003	40.596	-73.812	1	9.5	m	
R-EMAP Region 2 2003	2003	JB372	15-AUG-2003	40.596	-73.812	2	9.5	m	
R-EMAP Region 2 2003	2003	JB374	08-SEP-2003	40.624	-73.76	1	8.8	m	
R-EMAP Region 2 2003	2003	JB374	25-SEP-2003	40.624	-73.76	2	8.8	m	
R-EMAP Region 2 2003	2003	JB380	09-SEP-2003	40.629	-73.854	1	6.4	m	
R-EMAP Region 2 2003	2003	JB380	12-SEP-2003	40.629	-73.854	2	6.4	m	
R-EMAP Region 2 2003	2003	JB381	15-SEP-2003	40.601	-73.774	1	2.6	m	
R-EMAP Region 2 2003	2003	JB381	24-SEP-2003	40.601	-73.774	2	2.6	m	
R-EMAP Region 2 2003	2003	JB386	09-SEP-2003	40.604	-73.864	1	8.5	m	
R-EMAP Region 2 2003	2003	JB386	12-SEP-2003	40.604	-73.864	2	8.5	m	
R-EMAP Region 2 1993-94	1993	LS001	03-OCT-1993	41.056	-73.35	1	9.8	m	
R-EMAP Region 2 1993-94	1993	LS004	03-OCT-1993	41.015	-73.427	1	23.2	m	
R-EMAP Region 2 1993-94	1993	LS006	23-SEP-1993	41.081	-73.377	1	3.5	m	
R-EMAP Region 2 1993-94	1993	LS010	03-OCT-1993	40.979	-73.511	1	30.2	m	
R-EMAP Region 2 1993-94	1993	LS011	03-OCT-1993	40.972	-73.476	1	22.9	m	
R-EMAP Region 2 1993-94	1993	LS016	03-OCT-1993	40.948	-73.562	1	16.5	m	
R-EMAP Region 2 1993-94	1993	LS018	03-OCT-1993	40.947	-73.458	1	8.5	m	
R-EMAP Region 2 1993-94	1993	LS019	03-OCT-1993	40.919	-73.602	1	15.8	m	
R-EMAP Region 2 1993-94	1993	LS020	03-OCT-1993	40.911	-73.656	1	18.9	m	
R-EMAP Region 2 1993-94	1993	LS024	02-OCT-1993	41.018	-73.488	1	16.8	m	
R-EMAP Region 2 1993-94	1993	LS026	27-SEP-1993	41.002	-73.619	1	5.2	m	
R-EMAP Region 2 1993-94	1993	LS027	03-OCT-1993	40.982	-73.554	1	28.7	m	
R-EMAP Region 2 1993-94	1993	LS030	27-SEP-1993	40.95	-73.696	1	2.9	m	
R-EMAP Region 2 1993-94	1993	LS035	22-SEP-1993	40.833	-73.779	1	16.8	m	
R-EMAP Region 2 1993-94	1994	LS101	11-AUG-1994	41.05	-73.38	1	10.7	m	
R-EMAP Region 2 1993-94	1994	LS102	11-AUG-1994	41.022	-73.401	1	21.6	m	
R-EMAP Region 2 1993-94	1994	LS103	12-AUG-1994	41.006	-73.409	1	29.0	m	
R-EMAP Region 2 1993-94	1994	LS104	12-AUG-1994	40.99	-73.386	1	21.6	m	
R-EMAP Region 2 1993-94	1994	LS106	12-AUG-1994	40.972	-73.551	1	19.5	m	
R-EMAP Region 2 1993-94	1994	LS107	12-AUG-1994	40.966	-73.441	1	14.0	m	
R-EMAP Region 2 1993-94	1994	LS108	12-AUG-1994	40.957	-73.642	1	14.9	m	
R-EMAP Region 2 1993-94	1994	LS109	12-AUG-1994	40.949	-73.408	1	12.5	m	
R-EMAP Region 2 1993-94	1994	LS110	12-AUG-1994	40.934	-73.576	1	15.8	m	
R-EMAP Region 2 1993-94	1994	LS111	12-AUG-1994	40.917	-73.623	1	17.7	m	
R-EMAP Region 2 1993-94	1994	LS112	12-AUG-1994	40.91	-73.718	1	11.9	m	
R-EMAP Region 2 1993-94	1994	LS113	12-AUG-1994	40.869	-73.686	1	8.8	m	
R-EMAP Region 2 1993-94	1994	LS114	12-AUG-1994	40.85	-73.761	1	29.0	m	
R-EMAP Region 2 1993-94	1994	LS115	12-AUG-1994	40.95	-73.519	1	19.5	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2000	MA00-0009-C	23-AUG-2000	41.738	-70.622	1	6.0	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2000	MA00-0033-A	24-AUG-2000	41.442	-70.9	1	13.3	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2000	MA00-0035-B	13-SEP-2000	41.523	-71.065	1	6.1	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2000	MA00-0037-A	24-AUG-2000	41.513	-70.85	1	17.5	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2000	MA00-0039-A	13-SEP-2000	41.551	-71.061	1	1.5	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2000	MA00-0041-A	24-AUG-2000	41.584	-70.797	1	11.1	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2000	MA00-0045-A	24-AUG-2000	41.655	-70.745	1	5.3	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2000	MA00-0047-A	07-SEP-2000	41.734	-70.712	1	2.1	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2000	MA00-0049-A	18-SEP-2000	41.276	-70.207	1	0.5	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2000	MA00-0051-B	06-OCT-2000	41.36	-70.502	1	3.2	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2000	MA00-0053-A	22-SEP-2000	41.333	-70.028	1	2.3	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2000	MA00-0055-B	06-OCT-2000	41.433	-70.602	1	8.0	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2000	MA00-0057-C	29-SEP-2000	41.557	-70.526	1	2.2	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2000	MA00-0059-A	29-SEP-2000	41.613	-70.457	1	0.7	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2000	MA00-0061-C	29-SEP-2000	41.635	-70.242	1	1.0	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2000	MA00-0063-B	03-OCT-2000	41.72	-69.986	1	4.4	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2000	MA00-0069-A	25-JUL-2000	42.281	-70.883	1	2.0	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	MA00-0083-A	11-AUG-2000	41.732	-71.146	1	12.5	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	MA00-0085-A	15-AUG-2000	41.784	-71.118	1	3.5	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	MA00-0087-A	15-AUG-2000	41.815	-71.113	1	1.3	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	MA00-0089-B	15-AUG-2000	41.833	-71.109	1	3.0	m	
National Coastal Assessment-Northeast/Massachusetts Marine Fisheries	2000	MA00-0091-A	08-SEP-2000	42.45	-70.919	1	8.0	m	
National Coastal Assessment-Northeast/Massachusetts Marine Fisheries	2000	MA00-0093-A	08-SEP-2000	42.451	-70.911	1	11.0	m	
National Coastal Assessment-Northeast/Massachusetts Marine Fisheries	2000	MA00-0095-A	09-SEP-2000	42.698	-70.71	1	17.0	m	
National Coastal Assessment-Northeast/Massachusetts Marine Fisheries	2000	MA00-0097-A	09-SEP-2000	42.68	-70.707	1	8.0	m	
National Coastal Assessment-Northeast/Massachusetts Marine Fisheries	2000	MA00-0099-A	10-SEP-2000	42.026	-70.337	1	51.0	m	
National Coastal Assessment-Northeast/Massachusetts Marine Fisheries	2000	MA00-0101-A	10-SEP-2000	41.933	-70.38	1	38.0	m	
National Coastal Assessment-Northeast/Massachusetts Marine Fisheries	2000	MA00-0103-A	11-SEP-2000	41.79	-70.27	1	20.0	m	
National Coastal Assessment-Northeast/Massachusetts Marine Fisheries	2000	MA00-0105-A	11-SEP-2000	41.831	-70.123	1	13.0	m	
National Coastal Assessment-Northeast/Massachusetts Marine Fisheries	2000	MA00-0107-A	11-SEP-2000	41.9	-70.132	1	13.0	m	
National Coastal Assessment-Northeast/Massachusetts Marine Fisheries	2000	MA00-0109-A	11-SEP-2000	41.949	-70.095	1	9.0	m	
National Coastal Assessment-Northeast/Massachusetts Marine Fisheries	2000	MA00-0111-A	11-SEP-2000	41.879	-70.195	1	25.0	m	
National Coastal Assessment-Northeast/Massachusetts Marine Fisheries	2000	MA00-0113-A	12-SEP-2000	41.895	-70.414	1	32.0	m	
National Coastal Assessment-Northeast/Massachusetts Marine Fisheries	2000	MA00-0115-A	12-SEP-2000	41.896	-70.351	1	32.0	m	
National Coastal Assessment-Northeast/Massachusetts Marine Fisheries	2000	MA00-0117-A	12-SEP-2000	41.921	-70.273	1	34.0	m	
National Coastal Assessment-Northeast/Massachusetts Marine Fisheries	2000	MA00-0119-A	12-SEP-2000	41.949	-70.218	1	34.0	m	
National Coastal Assessment-Northeast/Massachusetts Marine Fisheries	2000	MA00-0121-A	12-SEP-2000	41.98	-70.138	1	27.0	m	
National Coastal Assessment-Northeast/Massachusetts Marine Fisheries	2000	MA00-0123-A	13-SEP-2000	41.994	-70.219	1	38.0	m	
National Coastal Assessment-Northeast/Massachusetts Marine Fisheries	2000	MA00-0125-A	20-SEP-2000	41.497	-70.849	1	17.0	m	
National Coastal Assessment-Northeast/Massachusetts Marine Fisheries	2000	MA00-0127-A	20-SEP-2000	41.539	-70.77	1	14.0	m	
National Coastal Assessment-Northeast/Massachusetts Marine Fisheries	2000	MA00-0129-A	20-SEP-2000	41.565	-70.676	1	15.0	m	
National Coastal Assessment-Northeast/Massachusetts Marine Fisheries	2000	MA00-0131-A	20-SEP-2000	41.657	-70.701	1	8.0	m	
National Coastal Assessment-Northeast/Massachusetts Marine Fisheries	2000	MA00-0133-A	20-SEP-2000	41.671	-70.729	1	6.0	m	
National Coastal Assessment-Northeast/Massachusetts Marine Fisheries	2000	MA00-0135-A	20-SEP-2000	41.593	-70.672	1	15.0	m	
National Coastal Assessment-Northeast/Massachusetts Marine Fisheries	2000	MA00-0137-A	06-SEP-2000	41.818	-70.525	1	10.0	m	
National Coastal Assessment-Northeast/Massachusetts Marine Fisheries	2000	MA00-0139-A	06-SEP-2000	41.845	-70.413	1	25.0	m	
National Coastal Assessment-Northeast/Massachusetts Marine Fisheries	2000	MA00-0141-A	06-SEP-2000	41.804	-70.386	1	21.0	m	
National Coastal Assessment-Northeast/Massachusetts Marine Fisheries	2000	MA00-0143-A	06-SEP-2000	41.748	-70.329	1	11.0	m	
National Coastal Assessment-Northeast/Massachusetts Marine Fisheries	2000	MA00-0145-A	06-SEP-2000	41.805	-70.491	1	18.0	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	MA01-0004-A	29-JUN-2001	42.551	-70.915	1	3.5	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	MA01-0010-A	23-JUL-2001	41.739	-70.616	1	8.5	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	MA01-0030-A	10-JUL-2001	42.032	-70.657	1	1.0	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	MA01-0034-C	21-AUG-2001	41.454	-70.807	1	4.7	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	MA01-0036-B	08-AUG-2001	41.479	-70.964	1	21.4	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	MA01-0038-A	08-AUG-2001	41.533	-70.695	1	10.8	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	MA01-0040-B	24-JUL-2001	41.642	-70.921	1	10.1	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	MA01-0042-A	24-JUL-2001	41.586	-70.686	1	13.2	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	MA01-0044-A	23-JUL-2001	41.653	-70.805	1	4.2	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	MA01-0046-B	23-JUL-2001	41.671	-70.636	1	7.2	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	MA01-0048-C	23-JUL-2001	41.709	-70.63	1	8.5	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	MA01-0050-A	28-SEP-2001	41.339	-70.773	1	1.4	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	MA01-0052-A	27-SEP-2001	41.298	-70.216	1	1.0	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	MA01-0054-A	27-SEP-2001	41.327	-70.003	1	1.8	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	MA01-0056-A	28-SEP-2001	41.449	-70.591	1	4.8	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	MA01-0058-B	30-SEP-2001	41.593	-70.459	1	1.2	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	MA01-0060-A	27-SEP-2001	41.641	-70.275	1	2.5	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	MA01-0062-B	04-OCT-2001	41.716	-69.975	1	4.1	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	MA01-0064-A	04-OCT-2001	41.748	-69.942	1	0.5	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	MA01-0068-A	05-JUL-2001	42.296	-71.043	1	8.2	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	MA01-0074-A	05-JUL-2001	42.433	-70.933	1	1.0	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	MA01-0076-A	27-JUN-2001	42.696	-70.805	1	2.0	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2001	MA01-0078-A	28-JUN-2001	42.664	-70.597	1	20.3	m	
National Coastal Assessment-Northeast/University of Rhode Island	2001	MA01-0082-A	02-AUG-2001	41.694	-71.189	1	10.5	m	
National Coastal Assessment-Northeast/University of Rhode Island	2001	MA01-0084-A	09-JUL-2001	41.725	-71.195	1	1.5	m	
National Coastal Assessment-Northeast/University of Rhode Island	2001	MA01-0088-A	10-JUL-2001	41.799	-71.119	1	1.3	m	
National Coastal Assessment-Northeast/University of Rhode Island	2001	MA01-0090-A	10-JUL-2001	41.875	-71.094	1	3.3	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2003	MA03-0051-B	09-SEP-2003	41.36	-70.502	1	2.8	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2003	MA03-0100-A	10-SEP-2003	41.331	-70.769	1	2.0	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2003	MA03-0103-C	18-AUG-2003	41.433	-70.953	1	12.0	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2003	MA03-0106-A	09-SEP-2003	41.336	-70.016	1	4.2	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2003	MA03-0109-A	18-AUG-2003	41.536	-70.724	1	15.2	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2003	MA03-0112-A	18-AUG-2003	41.552	-70.79	1	14.5	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2003	MA03-0115-A	01-OCT-2003	41.677	-70.917	1	1.5	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2003	MA03-0121-A	18-AUG-2003	41.736	-70.629	1	10.6	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2003	MA03-0130-A	24-SEP-2003	41.841	-69.951	1			
National Coastal Assessment-Northeast/University of Rhode Island	2003	MA03-0301-A	18-AUG-2003	41.713	-71.162	1	10.0	m	
National Coastal Assessment-Northeast/University of Rhode Island	2003	MA03-0306-B	09-SEP-2003	41.874	-71.093	1	3.3	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2004	MA04-0040-A	12-JUL-2004	41.643	-70.912	1	9.1	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2004	MA04-0101-A	03-SEP-2004	41.29	-70.224	1	2.5	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2004	MA04-0104-B	02-SEP-2004	41.352	-70.767	1	2.1	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2004	MA04-0107-A	02-SEP-2004	41.546	-71.062	1	1.2	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2004	MA04-0110-A	02-SEP-2004	41.459	-70.623	1	1.8	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2004	MA04-0113-A	12-JUL-2004	41.57	-70.721	1	11.0	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2004	MA04-0116-B	12-JUL-2004	41.654	-70.728	1	6.0	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2004	MA04-0119-B	08-SEP-2004	41.723	-69.935	1	0.1	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2004	MA04-0125-B	08-SEP-2004	41.732	-69.981	1			
National Coastal Assessment-Northeast/University of Rhode Island	2004	MA04-0300-A	15-JUL-2004	41.697	-71.184	1	12.4	m	
National Coastal Assessment-Northeast/University of Rhode Island	2004	MA04-0304-A	26-JUL-2004	41.778	-71.118	1	3.1	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2005	MA05-0001-A	26-AUG-2005	41.593	-70.716	1	11.8	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2005	MA05-0005-A	27-AUG-2005	41.513	-70.811	1	14.7	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2005	MA05-0007-A	26-AUG-2005	41.615	-70.89	1	3.9	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2005	MA05-0009-A	24-AUG-2005	41.698	-70.643	1	5.0	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2005	MA05-0013-A	27-AUG-2005	41.561	-70.705	1	13.5	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2005	MA05-0019-A	26-AUG-2005	41.64	-70.776	1	6.1	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2005	MA05-0020-A	27-AUG-2005	41.448	-70.902	1	11.0	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2006	MA06-0028-A	09-AUG-2006	41.678	-70.73	1	5.4	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2006	MA06-0029-A	09-AUG-2006	41.505	-70.862	1	16.4	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2006	MA06-0036-A	09-AUG-2006	41.516	-70.979	1	9.3	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2006	MA06-0042-A	09-AUG-2006	41.6	-70.645	1	9.0	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2006	MA06-0046-A	09-AUG-2006	41.566	-70.809	1	10.2	m	
National Coastal Assessment-Northeast/MA Coastal Zone Mgt/UMASS, Boston	2006	MA06-0050-A	09-AUG-2006	41.491	-70.843	1	15.0	m	
EMAP Mid-Atlantic Integrated Assessment/National Park Service	1997	MA97-0001	25-AUG-1997	38.327	-75.104	1	1.6	m	
EMAP Mid-Atlantic Integrated Assessment/National Park Service	1997	MA97-0003	26-AUG-1997	38.239	-75.209	1	1.3	m	
EMAP Mid-Atlantic Integrated Assessment/National Park Service	1997	MA97-0004	26-AUG-1997	38.253	-75.192	1	1.0	m	
EMAP Mid-Atlantic Integrated Assessment/National Park Service	1997	MA97-0005	27-AUG-1997	38.146	-75.286	1	0.8	m	
EMAP Mid-Atlantic Integrated Assessment/National Park Service	1997	MA97-0006	27-AUG-1997	38.105	-75.232	1	1.9	m	
EMAP Mid-Atlantic Integrated Assessment/National Park Service	1997	MA97-0007	05-SEP-1997	38.074	-75.361	1	1.0	m	
EMAP Mid-Atlantic Integrated Assessment/National Park Service	1997	MA97-0008	03-SEP-1997	37.981	-75.31	1	1.0	m	
EMAP Mid-Atlantic Integrated Assessment/National Park Service	1997	MA97-0009	02-SEP-1997	38.002	-75.385	1	2.0	m	
EMAP Mid-Atlantic Integrated Assessment/National Park Service	1997	MA97-0010	02-SEP-1997	37.984	-75.424	1	1.5	m	
EMAP Mid-Atlantic Integrated Assessment/National Park Service	1997	MA97-0011	28-AUG-1997	37.93	-75.391	1	3.6	m	
EMAP Mid-Atlantic Integrated Assessment/National Park Service	1997	MA97-0012	28-AUG-1997	37.915	-75.383	1	5.3	m	
EMAP Mid-Atlantic Integrated Assessment/National Park Service	1997	MA97-0013	29-AUG-1997	37.889	-75.372	1	2.8	m	
EMAP Mid-Atlantic Integrated Assessment/National Park Service	1997	MA97-0014	03-SEP-1997	38.067	-75.332	1	1.6	m	
EMAP Mid-Atlantic Integrated Assessment/National Park Service	1997	MA97-0015	08-SEP-1997	38.036	-75.268	1	1.8	m	
EMAP Mid-Atlantic Integrated Assessment/National Park Service	1997	MA97-0016	26-AUG-1997	38.215	-75.181	1	1.9	m	
EMAP Mid-Atlantic Integrated Assessment/National Park Service	1997	MA97-0017	25-AUG-1997	38.326	-75.1	1	2.6	m	
EMAP Mid-Atlantic Integrated Assessment/National Park Service	1997	MA97-0018	22-AUG-1997	38.285	-75.131	1	1.6	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0031	21-AUG-1997	38.206	-75.177	1	1.3	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0032	21-AUG-1997	38.228	-75.174	1	1.5	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0033	20-AUG-1997	38.246	-75.15	1	2.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0034	20-AUG-1997	38.264	-75.142	1	1.5	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0035	19-AUG-1997	38.282	-75.134	1	1.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0046	01-AUG-1997	37.375	-75.754	1	8.2	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0047	02-AUG-1997	37.703	-75.583	1	2.5	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0049	23-SEP-1997	37.931	-75.417	1	1.4	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0050	24-SEP-1997	37.876	-75.379	1	1.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0051	23-SEP-1997	37.908	-75.412	1	1.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0052	22-SEP-1997	37.956	-75.325	1	3.3	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0053	02-AUG-1997	37.305	-75.802	1	4.6	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0054	31-JUL-1997	37.173	-75.925	1	1.2	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0055	31-JUL-1997	37.214	-75.924	1	0.6	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0056	31-JUL-1997	37.333	-75.892	1	1.8	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0057	02-AUG-1997	37.623	-75.652	1	1.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0058	01-AUG-1997	37.458	-75.678	1	9.8	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0059	01-AUG-1997	37.367	-75.75	1	4.6	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0060	01-AUG-1997	37.399	-75.76	1	1.1	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0061	27-JUL-1997	37.294	-76.365	1	4.2	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0062	26-JUL-1997	37.304	-76.33	1	6.2	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0063	26-JUL-1997	37.331	-76.316	1	2.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0064	27-JUL-1997	37.321	-76.369	1	5.4	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0065	26-JUL-1997	37.333	-76.359	1	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0066	26-JUL-1997	37.341	-76.33	1	1.9	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0067	27-JUL-1997	37.336	-76.397	1	1.5	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0068	26-JUL-1997	37.348	-76.376	1	6.6	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0069	27-JUL-1997	37.368	-76.345	1	6.5	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0070	26-JUL-1997	37.365	-76.399	1	2.3	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0071	29-JUL-1997	37.312	-77.334	1	1.3	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0073	09-SEP-1997	38.568	-76.207	1	2.7	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0074	09-SEP-1997	38.745	-76.25	1	2.9	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0076	31-JUL-1997	37.303	-76.015	1	1.3	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0077	29-JUL-1997	37.301	-76.875	1	3.6	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0078	08-SEP-1997	38.929	-76.315	1	2.8	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0079	14-SEP-1997	39.507	-75.916	1	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0080	30-AUG-1997	37.482	-76.276	1	0.8	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0081	13-SEP-1997	37.848	-75.686	1	2.1	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0084	30-AUG-1997	37.644	-76.31	1	1.4	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0085	30-JUL-1997	36.887	-76.075	1	0.9	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0086	10-SEP-1997	38.115	-75.888	1	2.8	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0089	26-AUG-1997	39.214	-76.452	1	2.3	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0090	26-AUG-1997	39.248	-76.553	1	10.5	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0091	30-AUG-1997	37.522	-76.412	1	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0094	10-SEP-1997	38.346	-76.247	1	1.4	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0096	30-JUL-1997	37.083	-76.543	1	2.4	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0097	08-SEP-1997	38.877	-76.126	1	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0110	04-AUG-1997	39.08	-76.602	1	2.8	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0111	05-AUG-1997	39.074	-76.592	1	1.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0112	05-AUG-1997	39.063	-76.561	1	4.6	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0113	06-AUG-1997	39.059	-76.559	1	7.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0114	07-AUG-1997	39.059	-76.569	1	6.6	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0115	06-AUG-1997	39.057	-76.548	1	2.2	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0116	06-AUG-1997	39.052	-76.543	1	7.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0117	08-AUG-1997	39.048	-76.565	1	5.5	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0118	07-AUG-1997	39.047	-76.555	1	7.2	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0119	09-AUG-1997	39.048	-76.536	1	2.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0120	09-AUG-1997	39.043	-76.548	1	6.9	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0121	08-AUG-1997	39.043	-76.559	1	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0122	08-AUG-1997	39.035	-76.558	1	2.3	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0123	14-AUG-1997	39.034	-76.532	1	1.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0124	15-AUG-1997	39.034	-76.53	1	0.9	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0125	09-AUG-1997	39.034	-76.541	1	6.7	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0126	14-AUG-1997	39.03	-76.53	1	9.2	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0127	15-AUG-1997	39.022	-76.514	1	1.8	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0128	10-AUG-1997	39.017	-76.536	1	6.3	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0129	12-AUG-1997	39.013	-76.514	1	8.3	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0130	12-AUG-1997	39.007	-76.51	1	1.9	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0131	15-AUG-1997	39.004	-76.523	1	0.8	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0132	11-AUG-1997	39.003	-76.494	1	8.6	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0133	12-AUG-1997	38.998	-76.502	1	0.9	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0134	11-AUG-1997	38.989	-76.48	1	7.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0135	13-AUG-1997	38.977	-76.464	1	6.3	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0136	08-AUG-1997	38.974	-76.469	1	4.7	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0137	13-AUG-1997	38.969	-76.471	1	7.5	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0138	19-AUG-1997	38.967	-76.597	1	2.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0139	13-AUG-1997	38.962	-76.482	1	3.1	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0140	18-AUG-1997	38.956	-76.581	1	0.8	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0141	19-AUG-1997	38.956	-76.575	1	3.8	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0142	18-AUG-1997	38.953	-76.565	1	4.8	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0143	19-AUG-1997	38.952	-76.57	1	1.6	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0144	19-AUG-1997	38.951	-76.538	1	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0145	18-AUG-1997	38.95	-76.55	1	5.1	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0146	22-AUG-1997	38.949	-76.537	1	4.6	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0147	16-AUG-1997	38.941	-76.509	1	1.2	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0148	16-AUG-1997	38.939	-76.58	1	2.3	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0149	20-AUG-1997	38.938	-76.535	1	0.8	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0150	22-AUG-1997	38.933	-76.524	1	1.7	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0151	22-AUG-1997	38.932	-76.519	1	6.2	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0152	23-AUG-1997	38.929	-76.521	1	4.5	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0153	25-AUG-1997	38.926	-76.489	1	2.9	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0154	23-AUG-1997	38.925	-76.503	1	3.1	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0155	25-AUG-1997	38.923	-76.492	1	3.2	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0156	23-AUG-1997	38.918	-76.482	1	1.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0157	23-AUG-1997	38.915	-76.505	1	3.5	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0158	25-AUG-1997	38.913	-76.496	1	4.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0159	21-AUG-1997	38.912	-76.481	1	1.3	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0160	25-AUG-1997	38.91	-76.5	1	3.5	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0161	16-AUG-1997	38.909	-76.47	1	1.6	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0162	21-AUG-1997	38.907	-76.476	1	4.1	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0163	21-AUG-1997	38.903	-76.488	1	2.4	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0164	22-AUG-1997	38.899	-76.481	1	4.8	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0165	21-AUG-1997	38.893	-76.486	1	3.8	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0168	29-JUL-1997	37.571	-77.023	1	0.9	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0169	28-JUL-1997	37.569	-76.983	1	1.8	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0170	28-JUL-1997	37.567	-76.975	1	0.6	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0171	28-JUL-1997	37.566	-76.883	1	2.2	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0172	28-JUL-1997	37.563	-76.903	1	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0173	28-JUL-1997	37.561	-76.993	1	0.3	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0174	29-JUL-1997	37.56	-76.962	1	0.1	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0175	28-JUL-1997	37.559	-76.877	1	1.3	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0176	29-JUL-1997	37.549	-76.97	1	5.5	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0177	28-JUL-1997	37.548	-76.891	1	1.4	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0178	30-JUL-1997	37.547	-76.818	1	3.5	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0228	01-AUG-1997	37.319	-75.996	1	1.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0229	01-AUG-1997	37.318	-75.989	1	1.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0230	03-AUG-1997	37.316	-76.004	1	1.3	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0231	01-AUG-1997	37.314	-75.994	1	1.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0232	31-JUL-1997	37.312	-76.005	1	1.3	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0233	03-AUG-1997	37.306	-76.013	1	2.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0234	31-JUL-1997	37.303	-76.008	1	1.5	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0235	31-JUL-1997	37.3	-76.015	1	3.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0236	03-AUG-1997	37.291	-76.018	1	0.9	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0237	29-AUG-1997	38.147	-76.354	1	1.3	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0238	27-AUG-1997	38.139	-76.35	1	2.2	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0239	29-AUG-1997	38.131	-76.35	1	1.8	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0240	27-AUG-1997	38.125	-76.349	1	2.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0241	27-AUG-1997	38.121	-76.345	1	1.5	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0242	29-AUG-1997	38.12	-76.347	1	1.4	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0243	28-AUG-1997	38.115	-76.348	1	1.8	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0244	28-AUG-1997	38.116	-76.344	1	1.3	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0245	28-AUG-1997	38.115	-76.355	1	1.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0246	28-AUG-1997	38.113	-76.344	1	1.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0247	11-SEP-1997	38.189	-75.386	1	1.8	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0248	12-SEP-1997	38.186	-75.393	1	1.4	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0249	12-SEP-1997	38.145	-75.45	1	2.7	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0250	12-SEP-1997	38.143	-75.444	1	3.2	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0251	12-SEP-1997	38.054	-75.631	1	5.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0260	16-JUL-1997	39.545	-76.082	1	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0260	30-JUL-1997	39.545	-76.082	2	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0260	13-AUG-1997	39.545	-76.082	3	6.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0260	27-AUG-1997	39.545	-76.082	4	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0260	10-SEP-1997	39.545	-76.082	5	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0261	16-JUL-1997	39.44	-76.025	1	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0261	30-JUL-1997	39.44	-76.025	2	5.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0261	13-AUG-1997	39.44	-76.025	3	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0261	27-AUG-1997	39.44	-76.025	4	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0261	10-SEP-1997	39.44	-76.025	5	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0262	16-JUL-1997	39.347	-76.175	1	13.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0262	30-JUL-1997	39.347	-76.175	2	12.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0262	13-AUG-1997	39.347	-76.175	3	12.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0262	27-AUG-1997	39.347	-76.175	4	13.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0262	10-SEP-1997	39.347	-76.175	5	12.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0263	16-JUL-1997	39.248	-76.238	1	13.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0263	30-JUL-1997	39.248	-76.238	2	12.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0263	13-AUG-1997	39.248	-76.238	3	13.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0263	27-AUG-1997	39.248	-76.238	4	13.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0263	10-SEP-1997	39.248	-76.238	5	12.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0264	16-JUL-1997	39.163	-76.306	1	12.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0264	30-JUL-1997	39.163	-76.306	2	12.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0264	13-AUG-1997	39.163	-76.306	3	12.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0264	27-AUG-1997	39.163	-76.306	4	12.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0264	10-SEP-1997	39.163	-76.306	5	12.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0265	15-JUL-1997	39.003	-76.388	1	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0265	29-JUL-1997	39.003	-76.388	2	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0265	12-AUG-1997	39.003	-76.388	3	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0265	26-AUG-1997	39.003	-76.388	4	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0265	09-SEP-1997	39.003	-76.388	5	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0266	15-JUL-1997	39.002	-76.346	1	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0266	29-JUL-1997	39.002	-76.346	2	7.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0266	12-AUG-1997	39.002	-76.346	3	7.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0266	26-AUG-1997	39.002	-76.346	4	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0266	09-SEP-1997	39.002	-76.346	5	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0267	15-JUL-1997	38.995	-76.36	1	25.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0267	29-JUL-1997	38.995	-76.36	2	24.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0267	12-AUG-1997	38.995	-76.36	3	24.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0267	26-AUG-1997	38.995	-76.36	4	25.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0267	09-SEP-1997	38.995	-76.36	5	25.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0268	15-JUL-1997	38.825	-76.4	1	33.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0268	29-JUL-1997	38.825	-76.4	2	30.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0268	12-AUG-1997	38.825	-76.4	3	31.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0268	26-AUG-1997	38.825	-76.4	4	32.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0268	09-SEP-1997	38.825	-76.4	5	30.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0269	15-JUL-1997	38.816	-76.371	1	25.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0269	29-JUL-1997	38.816	-76.371	2	21.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0269	12-AUG-1997	38.816	-76.371	3	22.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0269	26-AUG-1997	38.816	-76.371	4	25.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0269	09-SEP-1997	38.816	-76.371	5	22.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0270	15-JUL-1997	38.813	-76.463	1	9.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0270	29-JUL-1997	38.813	-76.463	2	8.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0270	12-AUG-1997	38.813	-76.463	3	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0270	26-AUG-1997	38.813	-76.463	4	9.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0270	09-SEP-1997	38.813	-76.463	5	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0271	15-JUL-1997	38.645	-76.418	1	27.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0271	29-JUL-1997	38.645	-76.418	2	27.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0271	12-AUG-1997	38.645	-76.418	3	27.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0271	26-AUG-1997	38.645	-76.418	4	27.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0271	09-SEP-1997	38.645	-76.418	5	27.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0272	15-JUL-1997	38.645	-76.4	1	10.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0272	29-JUL-1997	38.645	-76.4	2	8.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0272	12-AUG-1997	38.645	-76.4	3	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0272	26-AUG-1997	38.645	-76.4	4	10.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0272	09-SEP-1997	38.645	-76.4	5	8.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0273	15-JUL-1997	38.643	-76.502	1	9.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0273	29-JUL-1997	38.643	-76.502	2	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0273	12-AUG-1997	38.643	-76.502	3	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0273	26-AUG-1997	38.643	-76.502	4	9.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0273	09-SEP-1997	38.643	-76.502	5	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0274	15-JUL-1997	38.556	-76.493	1	10.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0274	29-JUL-1997	38.556	-76.493	2	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0274	12-AUG-1997	38.556	-76.493	3	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0274	26-AUG-1997	38.556	-76.493	4	10.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0274	09-SEP-1997	38.556	-76.493	5	10.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0275	15-JUL-1997	38.556	-76.435	1	27.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0275	29-JUL-1997	38.556	-76.435	2	27.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0275	12-AUG-1997	38.556	-76.435	3	26.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0275	26-AUG-1997	38.556	-76.435	4	27.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0275	09-SEP-1997	38.556	-76.435	5	27.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0276	15-JUL-1997	38.556	-76.39	1	22.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0276	29-JUL-1997	38.556	-76.39	2	21.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0276	12-AUG-1997	38.556	-76.39	3	22.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0276	26-AUG-1997	38.556	-76.39	4	22.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0276	09-SEP-1997	38.556	-76.39	5	22.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0277	14-JUL-1997	38.413	-76.343	1	30.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0277	28-JUL-1997	38.413	-76.343	2	30.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0277	11-AUG-1997	38.413	-76.343	3	28.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0277	25-AUG-1997	38.413	-76.343	4	29.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0277	08-SEP-1997	38.413	-76.343	5	30.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0278	14-JUL-1997	38.318	-76.293	1	34.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0278	28-JUL-1997	38.318	-76.293	2	32.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0278	11-AUG-1997	38.318	-76.293	3	34.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0278	25-AUG-1997	38.318	-76.293	4	33.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0278	08-SEP-1997	38.318	-76.293	5	32.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0279	14-JUL-1997	38.137	-76.228	1	30.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0279	28-JUL-1997	38.137	-76.228	2	30.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0279	11-AUG-1997	38.137	-76.228	3	29.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0279	25-AUG-1997	38.137	-76.228	4	30.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0279	08-SEP-1997	38.137	-76.228	5	30.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0280	14-JUL-1997	38.021	-76.348	1	20.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0280	28-JUL-1997	38.021	-76.348	2	19.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0280	11-AUG-1997	38.021	-76.348	3	19.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0280	25-AUG-1997	38.021	-76.348	4	20.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0280	08-SEP-1997	38.021	-76.348	5	20.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0281	14-JUL-1997	37.912	-76.168	1	27.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0281	28-JUL-1997	37.912	-76.168	2	26.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0281	11-AUG-1997	37.912	-76.168	3	27.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0281	25-AUG-1997	37.912	-76.168	4	26.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0281	08-SEP-1997	37.912	-76.168	5	27.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0282	14-JUL-1997	37.908	-75.792	1	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0282	28-JUL-1997	37.908	-75.792	2	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0282	11-AUG-1997	37.908	-75.792	3	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0282	26-AUG-1997	37.908	-75.792	4	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0282	09-SEP-1997	37.908	-75.792	5	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0283	14-JUL-1997	37.813	-76.295	1	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0283	28-JUL-1997	37.813	-76.295	2	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0283	11-AUG-1997	37.813	-76.295	3	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0283	26-AUG-1997	37.813	-76.295	4	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0283	09-SEP-1997	37.813	-76.295	5	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0284	14-JUL-1997	37.8	-76.175	1	31.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0284	28-JUL-1997	37.8	-76.175	2	31.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0284	11-AUG-1997	37.8	-76.175	3	31.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0284	26-AUG-1997	37.8	-76.175	4	26.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0284	09-SEP-1997	37.8	-76.175	5	26.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0285	14-JUL-1997	37.793	-75.844	1	19.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0285	28-JUL-1997	37.793	-75.844	2	14.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0285	11-AUG-1997	37.793	-75.844	3	10.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0285	26-AUG-1997	37.793	-75.844	4	12.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0285	09-SEP-1997	37.793	-75.844	5	25.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0286	14-JUL-1997	37.692	-76.19	1	16.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0286	28-JUL-1997	37.692	-76.19	2	17.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0286	11-AUG-1997	37.692	-76.19	3	18.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0286	26-AUG-1997	37.692	-76.19	4	16.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0286	09-SEP-1997	37.692	-76.19	5	17.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0287	14-JUL-1997	37.683	-75.99	1	26.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0287	28-JUL-1997	37.683	-75.99	2	24.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0287	11-AUG-1997	37.683	-75.99	3	23.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0287	26-AUG-1997	37.683	-75.99	4	22.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0287	09-SEP-1997	37.683	-75.99	5	20.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0288	15-JUL-1997	37.597	-76.285	1	10.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0288	29-JUL-1997	37.597	-76.285	2	10.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0288	12-AUG-1997	37.597	-76.285	3	10.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0288	25-AUG-1997	37.597	-76.285	4	10.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0288	08-SEP-1997	37.597	-76.285	5	10.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0289	14-JUL-1997	37.775	-75.975	1	24.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0289	28-JUL-1997	37.775	-75.975	2	24.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0289	11-AUG-1997	37.775	-75.975	3	24.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0289	26-AUG-1997	37.775	-75.975	4	20.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0289	09-SEP-1997	37.775	-75.975	5	18.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0290	14-JUL-1997	37.581	-76.058	1	13.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0290	28-JUL-1997	37.581	-76.058	2	13.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0290	11-AUG-1997	37.581	-76.058	3	15.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0290	26-AUG-1997	37.581	-76.058	4	13.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0290	09-SEP-1997	37.581	-76.058	5	17.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0291	14-JUL-1997	37.531	-76.307	1	7.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0291	28-JUL-1997	37.531	-76.307	2	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0291	11-AUG-1997	37.531	-76.307	3	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0291	25-AUG-1997	37.531	-76.307	4	7.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0291	08-SEP-1997	37.531	-76.307	5	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0292	15-JUL-1997	37.487	-76.157	1	10.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0292	31-JUL-1997	37.487	-76.157	2	11.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0292	12-AUG-1997	37.487	-76.157	3	11.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0292	25-AUG-1997	37.487	-76.157	4	11.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0292	08-SEP-1997	37.487	-76.157	5	11.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0293	15-JUL-1997	37.411	-76.16	1	12.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0293	31-JUL-1997	37.411	-76.16	2	13.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0293	12-AUG-1997	37.411	-76.16	3	12.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0293	25-AUG-1997	37.411	-76.16	4	12.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0293	08-SEP-1997	37.411	-76.16	5	12.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0294	15-JUL-1997	37.411	-76.08	1	21.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0294	31-JUL-1997	37.411	-76.08	2	22.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0294	12-AUG-1997	37.411	-76.08	3	22.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0294	25-AUG-1997	37.411	-76.08	4	22.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0294	08-SEP-1997	37.411	-76.08	5	22.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0295	15-JUL-1997	37.411	-76.025	1	13.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0295	31-JUL-1997	37.411	-76.025	2	13.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0295	12-AUG-1997	37.411	-76.025	3	13.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0295	25-AUG-1997	37.411	-76.025	4	13.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0295	08-SEP-1997	37.411	-76.025	5	13.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0296	15-JUL-1997	37.312	-76.347	1	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0296	31-JUL-1997	37.312	-76.347	2	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0296	12-AUG-1997	37.312	-76.347	3	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0296	25-AUG-1997	37.312	-76.347	4	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0296	08-SEP-1997	37.312	-76.347	5	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0297	15-JUL-1997	37.242	-76.387	1	12.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0297	31-JUL-1997	37.242	-76.387	2	13.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0297	12-AUG-1997	37.242	-76.387	3	13.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0297	25-AUG-1997	37.242	-76.387	4	12.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0297	08-SEP-1997	37.242	-76.387	5	12.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0298	15-JUL-1997	37.236	-76.208	1	10.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0298	31-JUL-1997	37.236	-76.208	2	10.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0298	12-AUG-1997	37.236	-76.208	3	10.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0298	25-AUG-1997	37.236	-76.208	4	10.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0298	08-SEP-1997	37.236	-76.208	5	10.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0299	15-JUL-1997	37.229	-76.054	1	20.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0299	31-JUL-1997	37.229	-76.054	2	21.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0299	12-AUG-1997	37.229	-76.054	3	20.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0299	25-AUG-1997	37.229	-76.054	4	20.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0299	08-SEP-1997	37.229	-76.054	5	20.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0300	15-JUL-1997	37.177	-76.373	1	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0300	31-JUL-1997	37.177	-76.373	2	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0300	12-AUG-1997	37.177	-76.373	3	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0300	25-AUG-1997	37.177	-76.373	4	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0300	08-SEP-1997	37.177	-76.373	5	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0301	16-JUL-1997	37.117	-76.126	1	12.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0301	01-AUG-1997	37.117	-76.126	2	15.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0301	13-AUG-1997	37.117	-76.126	3	14.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0301	26-AUG-1997	37.117	-76.126	4	13.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0301	10-SEP-1997	37.117	-76.126	5	16.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0302	15-JUL-1997	37.11	-76.293	1	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0302	31-JUL-1997	37.11	-76.293	2	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0302	12-AUG-1997	37.11	-76.293	3	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0302	25-AUG-1997	37.11	-76.293	4	7.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0302	08-SEP-1997	37.11	-76.293	5	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0303	16-JUL-1997	37.058	-75.973	1	11.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0303	01-AUG-1997	37.058	-75.973	2	14.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0303	13-AUG-1997	37.058	-75.973	3	14.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0303	27-AUG-1997	37.058	-75.973	4	12.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0303	10-SEP-1997	37.058	-75.973	5	13.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0304	16-JUL-1997	36.997	-76.303	1	7.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0304	01-AUG-1997	36.997	-76.303	2	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0304	13-AUG-1997	36.997	-76.303	3	7.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0304	27-AUG-1997	36.997	-76.303	4	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0304	10-SEP-1997	36.997	-76.303	5	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0305	16-JUL-1997	36.993	-76.011	1	15.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0305	01-AUG-1997	36.993	-76.011	2	15.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0305	13-AUG-1997	36.993	-76.011	3	15.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0305	27-AUG-1997	36.993	-76.011	4	15.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0305	10-SEP-1997	36.993	-76.011	5	15.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0306	16-JUL-1997	36.988	-76.168	1	12.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0306	01-AUG-1997	36.988	-76.168	2	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0306	13-AUG-1997	36.988	-76.168	3	10.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0306	27-AUG-1997	36.988	-76.168	4	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0306	10-SEP-1997	36.988	-76.168	5	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0307	16-JUL-1997	36.945	-76.025	1	18.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0307	01-AUG-1997	36.945	-76.025	2	18.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0307	13-AUG-1997	36.945	-76.025	3	18.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0307	27-AUG-1997	36.945	-76.025	4	17.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0307	10-SEP-1997	36.945	-76.025	5	18.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0308	15-JUL-1997	37.588	-76.163	1	13.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0308	29-JUL-1997	37.588	-76.163	2	13.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0308	12-AUG-1997	37.588	-76.163	3	13.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0308	25-AUG-1997	37.588	-76.163	4	13.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0308	08-SEP-1997	37.588	-76.163	5	13.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0309	26-AUG-1997	39.589	-75.955	1	2.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0310	26-AUG-1997	39.548	-75.867	1	0.4	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0311	26-AUG-1997	39.533	-76.02	1	1.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0312	26-AUG-1997	39.531	-76.051	1	1.1	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0313	26-AUG-1997	39.526	-76.07	1	1.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0314	26-AUG-1997	39.514	-75.899	1	1.4	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0315	26-AUG-1997	39.455	-76.051	1	2.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0316	26-AUG-1997	39.449	-76.008	1	1.1	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0317	29-AUG-1997	39.444	-76.242	1	2.4	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0318	26-AUG-1997	39.437	-76.055	1	4.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0319	29-AUG-1997	39.419	-76.234	1	2.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0320	26-AUG-1997	39.408	-76.066	1	5.4	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0321	27-AUG-1997	39.376	-76.159	1	5.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0322	27-AUG-1997	39.36	-76.146	1	13.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0323	29-AUG-1997	39.346	-76.36	1	1.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0324	27-AUG-1997	39.349	-76.143	1	5.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0325	27-AUG-1997	39.321	-76.377	1	2.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0326	27-AUG-1997	39.317	-76.361	1	1.4	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0327	27-AUG-1997	39.308	-76.391	1	2.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0328	27-AUG-1997	39.292	-76.477	1	2.1	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0329	27-AUG-1997	39.28	-76.445	1	2.1	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0330	27-AUG-1997	39.245	-76.405	1	3.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0331	03-SEP-1997	39.241	-76.554	1	15.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0332	03-SEP-1997	39.205	-76.527	1	3.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0333	03-SEP-1997	39.198	-76.478	1	3.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0334	03-SEP-1997	39.193	-76.391	1	4.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0335	03-SEP-1997	39.194	-76.524	1	2.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0336	03-SEP-1997	39.184	-76.482	1	3.1	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0337	03-SEP-1997	39.18	-76.464	1	3.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0338	03-SEP-1997	39.178	-76.46	1	4.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0339	03-SEP-1997	39.177	-76.29	1	11.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0340	03-SEP-1997	39.172	-76.423	1	4.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0341	03-SEP-1997	39.172	-76.317	1	5.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0342	03-SEP-1997	39.155	-76.339	1	5.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0343	03-SEP-1997	39.152	-76.416	1	7.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0344	03-SEP-1997	39.111	-76.392	1	7.4	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0345	03-SEP-1997	39.091	-76.284	1	7.1	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0346	03-SEP-1997	39.089	-76.336	1	6.9	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0347	28-AUG-1997	39.086	-76.451	1	4.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0348	28-AUG-1997	39.083	-76.514	1	5.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0349	19-SEP-1997	39.084	-76.193	1	4.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0350	03-SEP-1997	39.08	-76.331	1	8.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0351	19-SEP-1997	39.076	-76.136	1	3.1	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0352	25-AUG-1997	39.057	-76.554	1	7.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0353	25-AUG-1997	39.055	-76.554	1	7.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0354	03-SEP-1997	39.051	-76.288	1	2.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0355	27-AUG-1997	39.241	-76.264	1	5.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0356	03-SEP-1997	39.046	-76.396	1	8.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0357	25-AUG-1997	39.041	-76.557	1	6.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0358	25-AUG-1997	39.036	-76.57	1	3.4	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0359	03-SEP-1997	39.032	-76.255	1	3.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0360	19-SEP-1997	39.015	-76.171	1	4.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0361	19-SEP-1997	39.009	-76.167	1	3.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0362	19-SEP-1997	39.185	-76.06	1	0.9	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0363	25-AUG-1997	39.0	-76.497	1	4.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0364	04-SEP-1997	38.921	-76.296	1	3.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0365	28-AUG-1997	38.917	-76.494	1	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0366	28-AUG-1997	38.912	-76.493	1	4.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0367	04-SEP-1997	38.906	-76.139	1	2.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0368	28-AUG-1997	38.893	-76.537	1	1.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0369	16-SEP-1997	38.254	-76.347	1	9.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0370	04-SEP-1997	38.846	-76.263	1	2.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0371	04-SEP-1997	38.837	-76.317	1	7.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0372	04-SEP-1997	38.829	-76.239	1	8.1	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0373	04-SEP-1997	38.823	-76.208	1	3.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0374	02-SEP-1997	38.722	-76.382	1	6.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0375	02-SEP-1997	38.713	-76.133	1	2.1	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0376	26-SEP-1997	38.701	-75.991	1	2.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0377	26-SEP-1997	38.691	-75.976	1	3.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0378	22-SEP-1997	38.675	-77.113	1	1.1	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0379	02-SEP-1997	38.678	-76.214	1	1.1	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0380	22-SEP-1997	38.646	-77.21	1	1.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0381	02-SEP-1997	38.649	-76.498	1	7.4	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0382	02-SEP-1997	38.608	-76.071	1	0.9	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0383	02-SEP-1997	38.604	-76.113	1	10.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0384	22-SEP-1997	38.584	-77.257	1	0.9	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0385	02-SEP-1997	38.592	-75.992	1	4.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0386	22-SEP-1997	38.568	-77.251	1	4.1	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0387	02-SEP-1997	38.577	-76.023	1	10.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0388	22-SEP-1997	38.553	-77.251	1	8.9	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0389	05-SEP-1997	38.379	-76.504	1	6.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0390	05-SEP-1997	38.547	-76.676	1	2.4	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0391	02-SEP-1997	38.534	-76.327	1	2.4	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0392	12-SEP-1997	38.507	-76.668	1	2.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0393	08-SEP-1997	38.49	-75.8	1	6.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0394	22-SEP-1997	38.467	-77.296	1	4.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0395	12-SEP-1997	38.476	-76.647	1	2.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0396	12-SEP-1997	38.462	-76.655	1	2.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0397	08-SEP-1997	38.469	-75.818	1	1.1	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0398	05-SEP-1997	38.46	-76.597	1	1.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0399	05-SEP-1997	38.457	-76.644	1	3.3	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0400	15-SEP-1997	39.964	-75.183	1	10.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0401	16-SEP-1997	39.953	-75.181	1	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0402	15-SEP-1997	39.946	-75.132	1	2.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0403	16-SEP-1997	39.944	-75.199	1	6.8	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0404	16-SEP-1997	39.932	-75.209	1	7.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0405	16-SEP-1997	39.922	-75.204	1	8.1	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0406	17-SEP-1997	39.911	-75.212	1	9.6	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0407	15-SEP-1997	39.907	-75.133	1	1.7	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0408	17-SEP-1997	39.895	-75.207	1	10.2	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0409	15-SEP-1997	39.892	-75.194	1	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0410	17-SEP-1997	39.893	-75.197	1	11.8	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1997	MA97-0411	15-SEP-1997	39.886	-75.196	1	10.8	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0412	16-SEP-1997	39.878	-75.15	1	4.6	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0413	16-SEP-1997	39.866	-75.203	1	3.7	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0414	16-SEP-1997	39.866	-75.208	1	5.6	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0415	17-SEP-1997	39.861	-75.299	1	2.6	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0416	12-SEP-1997	39.857	-75.244	1	13.7	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0417	16-SEP-1997	39.852	-75.268	1	8.5	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0418	16-SEP-1997	39.837	-75.351	1	5.7	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0419	12-SEP-1997	39.818	-75.384	1	14.9	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0420	12-SEP-1997	39.809	-75.403	1	14.0	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0421	12-SEP-1997	39.784	-75.435	1	2.0	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0422	12-SEP-1997	39.772	-75.478	1	2.0	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0423	12-SEP-1997	39.771	-75.458	1	4.3	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0424	12-SEP-1997	39.745	-75.492	1	11.0	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0425	11-SEP-1997	39.721	-75.489	1	4.0	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0426	11-SEP-1997	39.693	-75.511	1	6.4	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0427	10-SEP-1997	39.658	-75.549	1	7.0	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0428	11-SEP-1997	39.668	-75.547	1	4.9	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0429	18-SEP-1997	39.651	-75.48	1	0.5	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0430	18-SEP-1997	39.638	-75.482	1	0.7	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0431	18-SEP-1997	39.626	-75.48	1	0.6	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0432	18-SEP-1997	39.607	-75.465	1	1.9	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0433	18-SEP-1997	39.602	-75.477	1	1.5	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0434	06-OCT-1997	39.601	-75.589	1	2.7	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0435	06-OCT-1997	39.593	-75.59	1	4.6	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0436	18-SEP-1997	39.583	-75.479	1	2.5	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0437	19-SEP-1997	39.583	-75.49	1	0.6	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0438	19-SEP-1997	39.579	-75.497	1	1.0	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0439	19-SEP-1997	39.578	-75.482	1	1.9	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0440	06-OCT-1997	39.572	-75.535	1	3.1	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0441	19-SEP-1997	39.571	-75.503	1	2.6	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0442	06-OCT-1997	39.543	-75.564	1	4.0	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0443	06-OCT-1997	39.536	-75.531	1	3.4	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0444	08-OCT-1997	39.481	-75.584	1	1.8	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0445	08-OCT-1997	39.474	-75.544	1	4.6	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0446	10-SEP-1997	39.466	-75.564	1	10.1	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0447	23-SEP-1997	39.447	-75.506	1	1.5	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0448	23-SEP-1997	39.448	-75.571	1	1.2	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0449	10-SEP-1997	39.435	-75.542	1	11.6	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0450	07-OCT-1997	39.427	-75.475	1	4.9	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0452	07-OCT-1997	39.38	-75.435	1	6.1	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0453	07-OCT-1997	39.381	-75.518	1	0.4	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0454	09-SEP-1997	39.344	-75.485	1	2.7	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0455	08-SEP-1997	39.278	-75.365	1	12.2	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0456	09-SEP-1997	39.25	-75.288	1	6.7	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0457	23-SEP-1997	39.24	-75.424	1	2.4	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0458	09-SEP-1997	39.24	-75.234	1	5.9	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0459	09-SEP-1997	39.205	-75.224	1	4.4	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0460	09-SEP-1997	39.18	-75.354	1	4.0	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0461	08-SEP-1997	39.173	-75.268	1	14.3	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0462	08-SEP-1997	39.201	-75.108	1	1.9	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0463	06-SEP-1997	39.148	-75.017	1	4.6	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0464	09-SEP-1997	39.163	-75.35	1	4.0	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0465	08-SEP-1997	39.129	-75.252	1	7.0	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0466	06-SEP-1997	39.073	-75.038	1	4.5	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0467	06-SEP-1997	39.067	-74.991	1	5.8	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0468	06-SEP-1997	39.052	-75.069	1	8.2	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0469	08-SEP-1997	39.042	-75.227	1	8.5	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0470	06-SEP-1997	39.029	-75.014	1	4.7	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0471	05-SEP-1997	38.986	-75.036	1	12.2	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0472	05-SEP-1997	38.986	-75.298	1	2.1	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0473	02-SEP-1997	38.926	-74.814	1	4.5	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0474	08-SEP-1997	38.923	-75.124	1	16.5	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0475	05-SEP-1997	38.92	-75.21	1	4.6	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0476	02-SEP-1997	38.887	-74.9	1	4.4	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0477	02-SEP-1997	38.886	-74.94	1	4.3	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0478	05-SEP-1997	38.881	-75.031	1	10.1	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0479	05-SEP-1997	38.877	-75.137	1	19.5	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0480	02-SEP-1997	38.845	-75.001	1	4.9	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0481	05-SEP-1997	38.805	-75.117	1	9.2	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0482	05-SEP-1997	38.825	-75.077	1	19.5	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0483	03-SEP-1997	38.772	-75.046	1	18.9	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0484	02-SEP-1997	38.72	-75.068	1	10.1	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0485	03-SEP-1997	38.7	-75.029	1	12.8	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0486	03-SEP-1997	38.669	-75.06	1	7.3	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0487	04-SEP-1997	38.562	-75.042	1	10.7	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0488	04-SEP-1997	38.561	-75.004	1	12.2	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0489	04-SEP-1997	38.517	-75.033	1	14.0	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0490	15-SEP-1997	40.068	-74.911	1	2.0	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0491	15-SEP-1997	40.147	-74.723	1	3.7	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0492	15-SEP-1997	40.069	-74.91	1	1.1	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0493	15-SEP-1997	40.054	-74.975	1	3.3	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0494	15-SEP-1997	39.975	-75.085	1	5.8	m	
EMAP Mid-Atlantic Integrated Assessment/National Oceanic and Atmospheric Adm.	1997	MA97-0495	15-SEP-1997	40.027	-75.007	1	5.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0600	08-JUL-1997	38.918	-76.942	1			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0600	28-JUL-1997	38.918	-76.942	2			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0600	05-AUG-1997	38.918	-76.942	3			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0600	25-AUG-1997	38.918	-76.942	4			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0600	02-SEP-1997	38.918	-76.942	5			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0600	22-SEP-1997	38.918	-76.942	6			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0604	08-JUL-1997	38.909	-76.956	1			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0604	05-AUG-1997	38.909	-76.956	2			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0604	02-SEP-1997	38.909	-76.956	3			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0607	08-JUL-1997	38.899	-76.963	1			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0607	05-AUG-1997	38.899	-76.963	2			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0607	02-SEP-1997	38.899	-76.963	3			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0610	08-JUL-1997	38.884	-76.969	1			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0610	05-AUG-1997	38.884	-76.969	2			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0610	02-SEP-1997	38.884	-76.969	3			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0612	08-JUL-1997	38.877	-76.972	1			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0612	05-AUG-1997	38.877	-76.972	2			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0612	02-SEP-1997	38.877	-76.972	3			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0613	08-JUL-1997	38.877	-76.976	1			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0613	28-JUL-1997	38.877	-76.976	2			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0613	05-AUG-1997	38.877	-76.976	3			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0613	25-AUG-1997	38.877	-76.976	4			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0613	02-SEP-1997	38.877	-76.976	5			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0613	22-SEP-1997	38.877	-76.976	6			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0618	08-JUL-1997	38.87	-76.947	1			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0618	05-AUG-1997	38.87	-76.947	2			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0618	02-SEP-1997	38.87	-76.947	3			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0619	08-JUL-1997	38.853	-77.005	1			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0619	28-JUL-1997	38.853	-77.005	2			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0619	05-AUG-1997	38.853	-77.005	3			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0619	25-AUG-1997	38.853	-77.005	4			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0619	02-SEP-1997	38.853	-77.005	5			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0619	22-SEP-1997	38.853	-77.005	6			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0622	08-JUL-1997	38.861	-77.013	1			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0622	05-AUG-1997	38.861	-77.013	2			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0622	02-SEP-1997	38.861	-77.013	3			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0626	08-JUL-1997	38.851	-77.023	1			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0626	05-AUG-1997	38.851	-77.023	2			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0626	02-SEP-1997	38.851	-77.023	3			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0627	31-JUL-1997	39.283	-76.45	1	1.9	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0627	28-AUG-1997	39.283	-76.45	2	1.9	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0627	25-SEP-1997	39.283	-76.45	3	1.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0628	16-JUL-1997	38.058	-75.808	1	5.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0628	14-AUG-1997	38.058	-75.808	2	4.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0628	24-SEP-1997	38.058	-75.808	3	4.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0629	17-JUL-1997	39.467	-75.875	1	3.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0629	14-AUG-1997	39.467	-75.875	2	2.9	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0629	25-SEP-1997	39.467	-75.875	3	2.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0630	31-JUL-1997	39.433	-76.242	1	2.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0630	28-AUG-1997	39.433	-76.242	2	2.4	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0630	25-SEP-1997	39.433	-76.242	3	2.1	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0634	07-JUL-1997	38.325	-76.376	1	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0634	21-JUL-1997	38.325	-76.376	2	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0634	04-AUG-1997	38.325	-76.376	3	9.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0634	19-AUG-1997	38.325	-76.376	4	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0634	02-SEP-1997	38.325	-76.376	5	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0634	18-SEP-1997	38.325	-76.376	6	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0637	17-JUL-1997	39.258	-75.925	1	6.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0637	31-JUL-1997	39.258	-75.925	2	5.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0637	14-AUG-1997	39.258	-75.925	3	5.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0637	28-AUG-1997	39.258	-75.925	4	5.4	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0637	22-SEP-1997	39.258	-75.925	5	5.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0638	16-JUL-1997	38.992	-76.217	1	11.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0638	30-JUL-1997	38.992	-76.217	2	12.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0638	13-AUG-1997	38.992	-76.217	3	14.9	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0638	27-AUG-1997	38.992	-76.217	4	13.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0638	09-SEP-1997	38.992	-76.217	5	14.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0638	23-SEP-1997	38.992	-76.217	6	20.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0639	16-JUL-1997	38.971	-76.248	1	5.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0639	13-AUG-1997	38.971	-76.248	2	5.1	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0639	09-SEP-1997	38.971	-76.248	3	6.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0641	15-JUL-1997	37.312	-76.873	1	4.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0641	19-AUG-1997	37.312	-76.873	2	4.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0641	23-SEP-1997	37.312	-76.873	3	4.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0642	15-JUL-1997	38.65	-76.275	1	7.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0642	29-JUL-1997	38.65	-76.275	2	7.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0642	12-AUG-1997	38.65	-76.275	3	7.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0642	26-AUG-1997	38.65	-76.275	4	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0642	10-SEP-1997	38.65	-76.275	5	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0642	23-SEP-1997	38.65	-76.275	6	7.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0643	15-JUL-1997	38.533	-76.308	1	13.1	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0643	29-JUL-1997	38.533	-76.308	2	10.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0643	12-AUG-1997	38.533	-76.308	3	13.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0643	26-AUG-1997	38.533	-76.308	4	13.4	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0643	10-SEP-1997	38.533	-76.308	5	13.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0643	23-SEP-1997	38.533	-76.308	6	11.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0644	15-JUL-1997	38.583	-76.05	1	9.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0644	29-JUL-1997	38.583	-76.05	2	7.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0644	12-AUG-1997	38.583	-76.05	3	8.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0644	26-AUG-1997	38.583	-76.05	4	8.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0644	10-SEP-1997	38.583	-76.05	5	7.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0644	22-SEP-1997	38.583	-76.05	6	3.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0645	15-JUL-1997	38.567	-76.058	1	11.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0645	29-JUL-1997	38.567	-76.058	2	14.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0645	12-AUG-1997	38.567	-76.058	3	12.1	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0645	26-AUG-1997	38.567	-76.058	4	13.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0645	10-SEP-1997	38.567	-76.058	5	12.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0645	23-SEP-1997	38.567	-76.058	6	11.9	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0646	10-JUL-1997	37.693	-76.473	1	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0646	13-AUG-1997	37.693	-76.473	2	7.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0646	15-SEP-1997	37.693	-76.473	3	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0648	16-JUL-1997	38.883	-76.25	1	12.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0648	30-JUL-1997	38.883	-76.25	2	12.4	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0648	13-AUG-1997	38.883	-76.25	3	12.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0648	27-AUG-1997	38.883	-76.25	4	13.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0648	09-SEP-1997	38.883	-76.25	5	12.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0648	23-SEP-1997	38.883	-76.25	6	13.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0649	08-JUL-1997	36.841	-76.289	1	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0649	05-AUG-1997	36.841	-76.289	2	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0649	23-SEP-1997	36.841	-76.289	3	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0652	08-JUL-1997	36.882	-76.339	1	14.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0652	05-AUG-1997	36.882	-76.339	2	14.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0652	23-SEP-1997	36.882	-76.339	3	14.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0655	15-JUL-1997	36.903	-76.333	1	15.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0655	19-AUG-1997	36.903	-76.333	2	15.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0655	23-SEP-1997	36.903	-76.333	3	15.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0657	08-JUL-1997	36.813	-76.306	1	13.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0657	05-AUG-1997	36.813	-76.306	2	13.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0657	23-SEP-1997	36.813	-76.306	3	12.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0660	08-JUL-1997	36.77	-76.296	1	4.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0660	05-AUG-1997	36.77	-76.296	2	7.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0660	23-SEP-1997	36.77	-76.296	3	4.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0661	08-JUL-1997	36.843	-76.36	1	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0661	05-AUG-1997	36.843	-76.36	2	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0661	23-SEP-1997	36.843	-76.36	3	3.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0662	17-JUL-1997	39.525	-75.817	1	14.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0662	14-AUG-1997	39.525	-75.817	2	13.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0662	25-SEP-1997	39.525	-75.817	3	13.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0663	17-JUL-1997	39.508	-75.9	1	12.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0663	14-AUG-1997	39.508	-75.9	2	12.9	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0663	25-SEP-1997	39.508	-75.9	3	12.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0664	31-JUL-1997	39.383	-76.342	1	2.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0664	28-AUG-1997	39.383	-76.342	2	2.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0664	25-SEP-1997	39.383	-76.342	3	1.9	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0665	15-JUL-1997	37.207	-76.652	1	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0665	19-AUG-1997	37.207	-76.652	2	11.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0665	23-SEP-1997	37.207	-76.652	3	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0666	15-JUL-1997	37.058	-76.583	1	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0666	19-AUG-1997	37.058	-76.583	2	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0666	23-SEP-1997	37.058	-76.583	3	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0669	15-JUL-1997	36.99	-76.46	1	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0669	19-AUG-1997	36.99	-76.46	2	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0669	23-SEP-1997	36.99	-76.46	3	7.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0670	15-JUL-1997	36.955	-76.392	1	16.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0670	19-AUG-1997	36.955	-76.392	2	16.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0670	23-SEP-1997	36.955	-76.392	3	15.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0671	15-JUL-1997	37.21	-76.793	1	14.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0671	19-AUG-1997	37.21	-76.793	2	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0671	23-SEP-1997	37.21	-76.793	3	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0674	15-JUL-1997	37.531	-77.434	1			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0674	19-AUG-1997	37.531	-77.434	2			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0674	23-SEP-1997	37.531	-77.434	3			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0675	15-JUL-1997	37.45	-77.42	1	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0675	19-AUG-1997	37.45	-77.42	2	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0675	23-SEP-1997	37.45	-77.42	3	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0676	15-JUL-1997	37.403	-77.392	1	11.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0676	19-AUG-1997	37.403	-77.392	2	11.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0676	23-SEP-1997	37.403	-77.392	3	11.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0677	15-JUL-1997	37.311	-77.297	1	4.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0677	19-AUG-1997	37.311	-77.297	2	7.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0677	23-SEP-1997	37.311	-77.297	3	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0678	15-JUL-1997	37.313	-77.233	1	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0678	19-AUG-1997	37.313	-77.233	2	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0678	23-SEP-1997	37.313	-77.233	3	7.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0679	15-JUL-1997	37.3	-77.125	1	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0679	19-AUG-1997	37.3	-77.125	2	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0679	23-SEP-1997	37.3	-77.125	3	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0682	15-JUL-1997	37.275	-76.989	1	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0682	19-AUG-1997	37.275	-76.989	2	11.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0682	23-SEP-1997	37.275	-76.989	3	10.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0684	30-JUL-1997	39.075	-76.475	1	5.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0684	27-AUG-1997	39.075	-76.475	2	5.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0684	24-SEP-1997	39.075	-76.475	3	5.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0685	16-JUL-1997	38.142	-75.817	1	5.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0685	14-AUG-1997	38.142	-75.817	2	5.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0685	24-SEP-1997	38.142	-75.817	3	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0686	08-JUL-1997	37.723	-77.024	1	3.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0686	11-AUG-1997	37.723	-77.024	2	2.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0686	09-SEP-1997	37.723	-77.024	3	3.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0688	11-AUG-1997	37.572	-76.793	1	11.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0688	09-SEP-1997	37.572	-76.793	2	14.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0689	31-JUL-1997	39.3	-76.4	1	3.4	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0689	28-AUG-1997	39.3	-76.4	2	3.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0689	25-SEP-1997	39.3	-76.4	3	3.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0690	17-JUL-1997	38.533	-75.717	1	4.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0690	14-AUG-1997	38.533	-75.717	2	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0690	24-SEP-1997	38.533	-75.717	3	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0691	17-JUL-1997	38.333	-75.883	1	3.9	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0691	13-AUG-1997	38.333	-75.883	2	3.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0691	25-SEP-1997	38.333	-75.883	3	4.1	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0692	17-JUL-1997	39.575	-75.958	1	2.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0692	14-AUG-1997	39.575	-75.958	2	2.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0692	25-SEP-1997	39.575	-75.958	3	2.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0693	08-JUL-1997	37.525	-76.87	1	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0693	11-AUG-1997	37.525	-76.87	2	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0693	09-SEP-1997	37.525	-76.87	3			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0694	15-JUL-1997	39.208	-76.525	1	15.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0694	29-JUL-1997	39.208	-76.525	2	15.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0694	12-AUG-1997	39.208	-76.525	3	15.1	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0694	26-AUG-1997	39.208	-76.525	4	15.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0694	10-SEP-1997	39.208	-76.525	5	15.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0694	23-SEP-1997	39.208	-76.525	6	16.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0695	07-JUL-1997	38.425	-76.602	1	12.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0695	21-JUL-1997	38.425	-76.602	2	12.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0695	04-AUG-1997	38.425	-76.602	3	12.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0695	19-AUG-1997	38.425	-76.602	4	12.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0695	02-SEP-1997	38.425	-76.602	5	12.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0695	18-SEP-1997	38.425	-76.602	6	12.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0696	07-JUL-1997	38.379	-76.511	1	17.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0696	21-JUL-1997	38.379	-76.511	2	17.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0696	04-AUG-1997	38.379	-76.511	3	18.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0696	19-AUG-1997	38.379	-76.511	4	17.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0696	02-SEP-1997	38.379	-76.511	5	17.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0696	18-SEP-1997	38.379	-76.511	6	17.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0697	07-JUL-1997	38.341	-76.488	1	23.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0697	21-JUL-1997	38.341	-76.488	2	23.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0697	04-AUG-1997	38.341	-76.488	3	24.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0697	19-AUG-1997	38.341	-76.488	4	23.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0697	02-SEP-1997	38.341	-76.488	5	23.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0697	18-SEP-1997	38.341	-76.488	6	23.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0698	07-JUL-1997	38.312	-76.422	1	15.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0698	21-JUL-1997	38.312	-76.422	2	16.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0698	04-AUG-1997	38.312	-76.422	3	15.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0698	19-AUG-1997	38.312	-76.422	4	16.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0698	02-SEP-1997	38.312	-76.422	5	16.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0698	18-SEP-1997	38.312	-76.422	6	15.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0699	07-JUL-1997	38.491	-76.664	1	11.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0699	21-JUL-1997	38.491	-76.664	2	10.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0699	04-AUG-1997	38.491	-76.664	3	11.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0699	19-AUG-1997	38.491	-76.664	4	11.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0699	02-SEP-1997	38.491	-76.664	5	11.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0699	18-SEP-1997	38.491	-76.664	6	11.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0700	07-JUL-1997	38.81	-76.713	1			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0700	21-JUL-1997	38.81	-76.713	2			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0700	04-AUG-1997	38.81	-76.713	3			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0700	19-AUG-1997	38.81	-76.713	4			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0700	02-SEP-1997	38.81	-76.713	5			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0700	18-SEP-1997	38.81	-76.713	6			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0701	07-JUL-1997	38.773	-76.71	1	2.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0701	21-JUL-1997	38.773	-76.71	2	2.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0701	04-AUG-1997	38.773	-76.71	3			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0701	19-AUG-1997	38.773	-76.71	4			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0701	02-SEP-1997	38.773	-76.71	5			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0701	18-SEP-1997	38.773	-76.71	6	2.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0702	07-JUL-1997	38.71	-76.702	1	11.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0702	21-JUL-1997	38.71	-76.702	2	11.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0702	04-AUG-1997	38.71	-76.702	3	10.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0702	19-AUG-1997	38.71	-76.702	4	11.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0702	02-SEP-1997	38.71	-76.702	5	11.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0702	18-SEP-1997	38.71	-76.702	6	11.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0703	07-JUL-1997	38.658	-76.685	1	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0703	21-JUL-1997	38.658	-76.685	2	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0703	04-AUG-1997	38.658	-76.685	3	7.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0703	19-AUG-1997	38.658	-76.685	4	6.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0703	02-SEP-1997	38.658	-76.685	5	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0703	18-SEP-1997	38.658	-76.685	6	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0704	07-JUL-1997	38.582	-76.681	1	3.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0704	21-JUL-1997	38.582	-76.681	2	3.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0704	04-AUG-1997	38.582	-76.681	3	3.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0704	19-AUG-1997	38.582	-76.681	4	3.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0704	02-SEP-1997	38.582	-76.681	5	3.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0704	18-SEP-1997	38.582	-76.681	6	3.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0705	07-JUL-1997	38.785	-76.714	1	1.1	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0705	21-JUL-1997	38.785	-76.714	2	1.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0705	04-AUG-1997	38.785	-76.714	3			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0705	19-AUG-1997	38.785	-76.714	4			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0705	02-SEP-1997	38.785	-76.714	5			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0705	18-SEP-1997	38.785	-76.714	6	1.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0707	17-JUL-1997	38.083	-75.567	1	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0707	14-AUG-1997	38.083	-75.567	2	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0707	24-SEP-1997	38.083	-75.567	3	4.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0708	16-JUL-1997	37.942	-75.767	1	4.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0708	31-JUL-1997	37.942	-75.767	2	3.9	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0708	14-AUG-1997	37.942	-75.767	3	4.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0708	28-AUG-1997	37.942	-75.767	4	4.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0708	10-SEP-1997	37.942	-75.767	5	4.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0708	24-SEP-1997	37.942	-75.767	6	3.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0709	14-JUL-1997	38.167	-76.583	1	12.4	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0709	28-JUL-1997	38.167	-76.583	2	11.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0709	11-AUG-1997	38.167	-76.583	3	12.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0709	25-AUG-1997	38.167	-76.583	4	12.4	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0709	09-SEP-1997	38.167	-76.583	5	12.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0709	22-SEP-1997	38.167	-76.583	6	12.9	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0710	14-JUL-1997	38.565	-77.194	1	7.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0710	28-JUL-1997	38.565	-77.194	2	7.4	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0710	11-AUG-1997	38.565	-77.194	3	6.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0710	25-AUG-1997	38.565	-77.194	4	6.1	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0710	08-SEP-1997	38.565	-77.194	5	7.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0710	22-SEP-1997	38.565	-77.194	6	6.9	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0711	14-JUL-1997	38.588	-77.119	1			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0711	28-JUL-1997	38.588	-77.119	2			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0711	11-AUG-1997	38.588	-77.119	3			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0711	25-AUG-1997	38.588	-77.119	4			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0711	08-SEP-1997	38.588	-77.119	5			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0711	22-SEP-1997	38.588	-77.119	6			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0722	14-JUL-1997	38.698	-76.987	1			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0722	28-JUL-1997	38.698	-76.987	2			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0722	11-AUG-1997	38.698	-76.987	3			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0722	25-AUG-1997	38.698	-76.987	4			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0722	08-SEP-1997	38.698	-76.987	5			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0722	22-SEP-1997	38.698	-76.987	6			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0723	14-JUL-1997	38.918	-77.105	1			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0723	11-AUG-1997	38.918	-77.105	2			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0723	08-SEP-1997	38.918	-77.105	3			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0731	14-JUL-1997	38.902	-77.07	1			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0731	28-JUL-1997	38.902	-77.07	2			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0731	11-AUG-1997	38.902	-77.07	3			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0731	25-AUG-1997	38.902	-77.07	4			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0731	08-SEP-1997	38.902	-77.07	5			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0731	22-SEP-1997	38.902	-77.07	6			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0742	14-JUL-1997	38.874	-77.043	1			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0742	28-JUL-1997	38.874	-77.043	2			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0742	11-AUG-1997	38.874	-77.043	3			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0742	25-AUG-1997	38.874	-77.043	4			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0742	08-SEP-1997	38.874	-77.043	5			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0742	22-SEP-1997	38.874	-77.043	6			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0750	14-JUL-1997	38.85	-77.023	1			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0750	28-JUL-1997	38.85	-77.023	2			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0750	11-AUG-1997	38.85	-77.023	3			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0750	25-AUG-1997	38.85	-77.023	4			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0750	08-SEP-1997	38.85	-77.023	5			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0750	22-SEP-1997	38.85	-77.023	6			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0758	14-JUL-1997	38.822	-77.031	1			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0758	11-AUG-1997	38.822	-77.031	2			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0758	08-SEP-1997	38.822	-77.031	3			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0765	14-JUL-1997	38.795	-77.037	1			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0765	11-AUG-1997	38.795	-77.037	2			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0765	08-SEP-1997	38.795	-77.037	3			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0772	14-JUL-1997	38.77	-77.032	1			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0772	11-AUG-1997	38.77	-77.032	2			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0772	08-SEP-1997	38.77	-77.032	3			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0773	07-JUL-1997	38.887	-77.04	1			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0773	04-AUG-1997	38.887	-77.04	2			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0773	09-SEP-1997	38.887	-77.04	3			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0777	08-JUL-1997	38.874	-77.023	1			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0777	05-AUG-1997	38.874	-77.023	2			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0777	02-SEP-1997	38.874	-77.023	3			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0782	14-JUL-1997	38.403	-77.269	1	7.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0782	28-JUL-1997	38.403	-77.269	2	7.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0782	11-AUG-1997	38.403	-77.269	3	7.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0782	25-AUG-1997	38.403	-77.269	4	6.9	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0782	08-SEP-1997	38.403	-77.269	5	7.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0782	22-SEP-1997	38.403	-77.269	6	7.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0783	14-JUL-1997	38.352	-77.205	1	9.1	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0783	28-JUL-1997	38.352	-77.205	2	9.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0783	11-AUG-1997	38.352	-77.205	3	10.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0783	25-AUG-1997	38.352	-77.205	4	9.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0783	08-SEP-1997	38.352	-77.205	5	10.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0783	22-SEP-1997	38.352	-77.205	6	9.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0785	14-JUL-1997	38.363	-76.991	1	14.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0785	28-JUL-1997	38.363	-76.991	2	15.4	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0785	11-AUG-1997	38.363	-76.991	3	14.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0785	25-AUG-1997	38.363	-76.991	4	14.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0785	08-SEP-1997	38.363	-76.991	5	15.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0785	22-SEP-1997	38.363	-76.991	6	15.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0787	14-JUL-1997	38.706	-77.049	1	18.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0787	28-JUL-1997	38.706	-77.049	2	19.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0787	11-AUG-1997	38.706	-77.049	3	19.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0787	25-AUG-1997	38.706	-77.049	4	18.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0787	08-SEP-1997	38.706	-77.049	5	20.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0787	22-SEP-1997	38.706	-77.049	6	18.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0788	14-JUL-1997	38.691	-77.111	1	8.1	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0788	28-JUL-1997	38.691	-77.111	2	7.9	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0788	11-AUG-1997	38.691	-77.111	3	8.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0788	25-AUG-1997	38.691	-77.111	4	8.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0788	08-SEP-1997	38.691	-77.111	5	8.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0788	22-SEP-1997	38.691	-77.111	6	8.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0789	14-JUL-1997	38.608	-77.174	1	11.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0789	28-JUL-1997	38.608	-77.174	2	11.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0789	11-AUG-1997	38.608	-77.174	3	12.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0789	25-AUG-1997	38.608	-77.174	4	12.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0789	08-SEP-1997	38.608	-77.174	5	12.9	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0789	22-SEP-1997	38.608	-77.174	6	12.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0790	14-JUL-1997	38.53	-77.266	1	8.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0790	28-JUL-1997	38.53	-77.266	2	8.4	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0790	11-AUG-1997	38.53	-77.266	3	8.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0790	25-AUG-1997	38.53	-77.266	4	8.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0790	08-SEP-1997	38.53	-77.266	5	8.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0790	22-SEP-1997	38.53	-77.266	6	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0792	10-JUL-1997	37.761	-76.621	1	7.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0792	13-AUG-1997	37.761	-76.621	2	7.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0792	15-SEP-1997	37.761	-76.621	3	7.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0793	10-JUL-1997	37.67	-76.554	1	14.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0793	13-AUG-1997	37.67	-76.554	2	15.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0793	15-SEP-1997	37.67	-76.554	3	14.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0796	10-JUL-1997	37.633	-76.463	1	11.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0796	13-AUG-1997	37.633	-76.463	2	11.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0796	15-SEP-1997	37.633	-76.463	3	11.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0799	10-JUL-1997	37.92	-76.822	1	4.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0799	13-AUG-1997	37.92	-76.822	2	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0799	10-SEP-1997	37.92	-76.822	3	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0802	10-JUL-1997	37.808	-76.713	1	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0802	13-AUG-1997	37.808	-76.713	2	4.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0802	10-SEP-1997	37.808	-76.713	3	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0805	10-JUL-1997	38.246	-77.234	1	3.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0805	18-AUG-1997	38.246	-77.234	2	3.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0805	15-SEP-1997	38.246	-77.234	3	3.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0808	10-JUL-1997	38.245	-77.326	1	3.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0808	18-AUG-1997	38.245	-77.326	2	3.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0808	15-SEP-1997	38.245	-77.326	3	3.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0809	10-JUL-1997	38.175	-77.189	1	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0809	18-AUG-1997	38.175	-77.189	2	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0809	15-SEP-1997	38.175	-77.189	3	4.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0810	10-JUL-1997	38.112	-77.052	1	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0810	13-AUG-1997	38.112	-77.052	2	4.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0810	10-SEP-1997	38.112	-77.052	3	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0811	10-JUL-1997	38.019	-76.908	1	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0811	13-AUG-1997	38.019	-76.908	2	7.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0811	10-SEP-1997	38.019	-76.908	3	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0812	30-JUL-1997	38.883	-76.533	1	2.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0812	27-AUG-1997	38.883	-76.533	2	2.9	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0812	24-SEP-1997	38.883	-76.533	3	2.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0813	30-JUL-1997	38.85	-76.533	1	3.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0813	27-AUG-1997	38.85	-76.533	2	3.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0813	24-SEP-1997	38.85	-76.533	3	3.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0814	07-JUL-1997	38.986	-77.064	1			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0814	04-AUG-1997	38.986	-77.064	2			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0814	09-SEP-1997	38.986	-77.064	3			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0817	07-JUL-1997	38.928	-77.05	1			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0817	04-AUG-1997	38.928	-77.05	2			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0817	09-SEP-1997	38.928	-77.05	3			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0818	31-JUL-1997	39.367	-75.883	1	6.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0818	28-AUG-1997	39.367	-75.883	2	6.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0818	24-SEP-1997	39.367	-75.883	3	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0819	08-JUL-1997	39.659	-76.174	1			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0819	05-AUG-1997	39.659	-76.174	2			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0819	15-SEP-1997	39.659	-76.174	3			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0820	17-JUL-1997	38.283	-76.017	1	7.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0820	13-AUG-1997	38.283	-76.017	2	7.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0820	25-SEP-1997	38.283	-76.017	3	7.1	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0821	17-JUL-1997	38.2	-75.975	1	13.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0821	31-JUL-1997	38.2	-75.975	2	13.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0821	13-AUG-1997	38.2	-75.975	3	14.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0821	28-AUG-1997	38.2	-75.975	4	14.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0821	10-SEP-1997	38.2	-75.975	5	14.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0821	25-SEP-1997	38.2	-75.975	6	13.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0822	16-JUL-1997	37.967	-75.933	1	27.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0822	31-JUL-1997	37.967	-75.933	2	29.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0822	14-AUG-1997	37.967	-75.933	3	28.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0822	28-AUG-1997	37.967	-75.933	4	28.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0822	10-SEP-1997	37.967	-75.933	5	27.9	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0822	24-SEP-1997	37.967	-75.933	6	26.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0823	17-JUL-1997	38.267	-75.792	1	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0823	13-AUG-1997	38.267	-75.792	2	8.1	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0823	25-SEP-1997	38.267	-75.792	3	8.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0824	08-JUL-1997	37.418	-76.693	1	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0824	11-AUG-1997	37.418	-76.693	2	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0824	09-SEP-1997	37.418	-76.693	3			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0825	08-JUL-1997	37.292	-76.558	1	12.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0825	11-AUG-1997	37.292	-76.558	2	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0825	09-SEP-1997	37.292	-76.558	3			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0828	08-JUL-1997	37.235	-76.485	1	15.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0828	11-AUG-1997	37.235	-76.485	2	20.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0828	09-SEP-1997	37.235	-76.485	3			
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0831	08-JUL-1997	37.58	-77.022	1	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0831	11-AUG-1997	37.58	-77.022	2	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0831	09-SEP-1997	37.58	-77.022	3	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0833	08-JUL-1997	37.507	-76.788	1	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0833	11-AUG-1997	37.507	-76.788	2	3.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0833	09-SEP-1997	37.507	-76.788	3	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0835	05-SEP-1997	38.451	-76.631	1	4.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0836	05-SEP-1997	38.445	-76.607	1	2.1	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0837	05-SEP-1997	38.437	-76.619	1	5.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0838	05-SEP-1997	38.409	-76.544	1	2.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0839	05-SEP-1997	38.406	-76.567	1	5.9	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0840	05-SEP-1997	38.404	-76.564	1	6.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0841	05-SEP-1997	38.394	-76.539	1	8.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0842	05-SEP-1997	38.393	-76.561	1	2.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0843	05-SEP-1997	38.391	-76.521	1	6.4	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0844	26-SEP-1997	38.379	-76.881	1	1.4	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0845	05-SEP-1997	38.37	-76.473	1	1.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0846	22-SEP-1997	38.355	-77.221	1	7.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0847	22-SEP-1997	38.342	-77.259	1	3.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0848	08-SEP-1997	38.361	-75.86	1	3.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0849	05-SEP-1997	38.347	-76.504	1	2.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0850	05-SEP-1997	38.343	-76.476	1	7.9	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0851	08-SEP-1997	38.342	-75.875	1	2.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0852	05-SEP-1997	38.419	-76.56	1	2.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0853	08-SEP-1997	38.333	-75.88	1	1.4	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0854	04-SEP-1997	38.319	-76.424	1	7.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0855	26-SEP-1997	38.306	-76.831	1	4.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0856	05-SEP-1997	38.376	-76.516	1	7.9	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0857	04-SEP-1997	38.303	-76.462	1	2.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0858	08-SEP-1997	38.305	-76.046	1	1.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0859	04-SEP-1997	38.299	-76.434	1	8.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0860	04-SEP-1997	38.297	-76.448	1	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0861	17-SEP-1997	38.259	-75.824	1	1.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0862	17-SEP-1997	38.239	-75.864	1	2.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0863	16-SEP-1997	38.227	-76.348	1	9.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0864	16-SEP-1997	38.219	-76.846	1	6.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0865	17-SEP-1997	38.201	-76.017	1	2.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0866	16-SEP-1997	38.19	-76.827	1	6.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0867	16-SEP-1997	38.186	-76.811	1	6.9	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0868	16-SEP-1997	38.187	-76.759	1	8.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0869	16-SEP-1997	38.182	-76.71	1	7.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0870	16-SEP-1997	38.173	-76.552	1	5.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0871	16-SEP-1997	38.166	-76.745	1	2.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0872	17-SEP-1997	38.168	-76.001	1	2.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0873	17-SEP-1997	38.148	-77.083	1	6.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0874	17-SEP-1997	38.151	-76.121	1	5.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0875	17-SEP-1997	38.13	-75.841	1	1.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0876	17-SEP-1997	38.128	-75.841	1	1.4	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0877	15-SEP-1997	38.102	-76.57	1	7.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0878	17-SEP-1997	38.09	-76.082	1	1.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0879	02-SEP-1997	38.621	-76.222	1	1.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0880	16-SEP-1997	38.225	-76.706	1	5.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0881	17-SEP-1997	38.065	-75.896	1	7.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0882	15-SEP-1997	38.058	-76.483	1	11.2	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0883	15-SEP-1997	38.053	-76.49	1	9.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0884	15-SEP-1997	38.052	-76.457	1	11.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0885	17-SEP-1997	38.048	-76.176	1	5.9	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0886	17-SEP-1997	38.049	-75.813	1	1.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0887	17-SEP-1997	38.045	-75.844	1	2.1	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0888	17-SEP-1997	38.022	-76.181	1	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0889	15-SEP-1997	38.015	-76.439	1	6.9	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0890	17-SEP-1997	38.008	-76.137	1	5.1	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0891	15-SEP-1997	38.003	-76.282	1	11.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0892	17-SEP-1997	37.99	-76.902	1	3.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0893	17-SEP-1997	37.975	-75.978	1	1.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0894	15-SEP-1997	37.964	-76.388	1	3.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0895	15-SEP-1997	37.96	-76.291	1	11.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0896	17-SEP-1997	37.944	-76.857	1	3.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0897	17-SEP-1997	37.941	-76.849	1	3.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0898	17-SEP-1997	37.917	-76.829	1	1.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0899	12-AUG-1997	37.915	-76.151	1	21.9	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0900	12-AUG-1997	37.872	-76.19	1	9.4	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0901	04-AUG-1997	37.209	-76.344	1	7.9	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0902	17-SEP-1997	37.867	-76.767	1	7.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0903	12-AUG-1997	37.849	-76.01	1	2.4	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0904	18-SEP-1997	37.839	-76.736	1	3.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0905	18-SEP-1997	37.823	-76.731	1	4.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0906	18-SEP-1997	37.808	-76.712	1	5.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0907	18-SEP-1997	37.804	-76.693	1	6.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0908	18-SEP-1997	37.795	-76.701	1	3.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0909	12-AUG-1997	37.782	-76.171	1	22.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0910	28-AUG-1997	37.776	-76.626	1	4.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0911	28-AUG-1997	37.758	-76.649	1	4.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0912	28-AUG-1997	37.748	-76.604	1	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0913	28-AUG-1997	37.724	-76.59	1	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0914	28-AUG-1997	37.715	-76.557	1	3.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0915	28-AUG-1997	37.694	-76.573	1	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0916	16-SEP-1997	37.687	-76.917	1	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0917	28-AUG-1997	37.678	-76.556	1	11.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0918	11-AUG-1997	37.681	-75.927	1	5.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0919	28-AUG-1997	37.656	-76.477	1	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0920	12-AUG-1997	37.659	-76.092	1	11.9	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0921	11-AUG-1997	37.646	-76.051	1	13.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0922	28-AUG-1997	37.633	-76.42	1	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0923	28-AUG-1997	37.632	-76.455	1	23.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0924	28-AUG-1997	37.626	-76.522	1	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0925	28-AUG-1997	37.622	-76.46	1	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0926	28-AUG-1997	37.61	-76.41	1	9.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0927	28-AUG-1997	37.592	-76.367	1	12.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0928	11-AUG-1997	37.591	-76.049	1	14.9	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0929	16-SEP-1997	37.558	-76.876	1	2.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0930	16-SEP-1997	37.556	-76.86	1	5.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0931	16-SEP-1997	37.538	-76.945	1	7.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0932	11-AUG-1997	37.52	-76.271	1	5.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0933	11-AUG-1997	37.519	-76.159	1	11.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0934	16-SEP-1997	37.5	-76.78	1	4.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0935	16-SEP-1997	37.499	-76.779	1	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0936	11-AUG-1997	37.493	-76.183	1	10.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0937	26-AUG-1997	37.433	-76.726	1	3.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0938	11-AUG-1997	37.427	-76.091	1	27.1	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0939	26-AUG-1997	37.397	-76.661	1	3.4	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0940	11-AUG-1997	37.402	-76.03	1	13.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0941	04-AUG-1997	37.395	-76.217	1	3.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0942	26-AUG-1997	37.38	-76.673	1	3.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0943	26-AUG-1997	37.38	-76.673	1	3.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0944	11-AUG-1997	37.378	-76.026	1	10.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0945	26-AUG-1997	37.369	-76.644	1	3.4	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0946	16-SEP-1997	37.526	-76.803	1	4.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0947	04-AUG-1997	37.366	-76.232	1	8.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0948	04-AUG-1997	37.346	-76.206	1	8.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0949	26-AUG-1997	37.341	-76.603	1	3.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0950	26-AUG-1997	37.456	-76.74	1	3.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0951	21-AUG-1997	37.316	-77.223	1	2.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0952	26-AUG-1997	37.312	-76.615	1	2.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0953	26-AUG-1997	37.307	-76.586	1	6.1	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0954	04-AUG-1997	37.146	-76.182	1	11.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0955	04-AUG-1997	37.3	-76.302	1	5.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0956	26-AUG-1997	37.277	-76.575	1	1.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0957	04-AUG-1997	37.282	-76.061	1	9.1	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0958	26-AUG-1997	37.276	-76.541	1	16.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0959	04-AUG-1997	37.276	-76.322	1	4.9	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0960	26-AUG-1997	37.257	-76.529	1	13.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0961	26-AUG-1997	37.254	-76.525	1	13.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0962	26-AUG-1997	37.253	-76.514	1	10.4	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0963	26-AUG-1997	37.246	-76.487	1	3.9	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0964	26-AUG-1997	37.245	-76.503	1	3.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0965	21-AUG-1997	37.238	-76.902	1	2.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0966	21-AUG-1997	37.232	-76.809	1	3.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0967	26-AUG-1997	37.234	-76.456	1	14.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0968	21-AUG-1997	37.217	-76.917	1	7.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0969	26-AUG-1997	37.224	-76.453	1	1.9	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0970	11-AUG-1997	37.225	-76.111	1	12.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0971	21-AUG-1997	37.212	-76.907	1	1.1	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0972	21-AUG-1997	37.209	-76.714	1	2.5	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0973	21-AUG-1997	37.184	-76.739	1	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0974	09-SEP-1997	37.181	-76.622	1	2.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0975	09-SEP-1997	37.148	-76.621	1	2.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0976	04-AUG-1997	37.143	-76.196	1	11.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0977	11-AUG-1997	37.132	-76.037	1	7.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0978	09-SEP-1997	37.106	-76.642	1	4.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0979	09-SEP-1997	37.078	-76.634	1	5.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0980	25-AUG-1997	36.96	-76.475	1	1.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0981	25-AUG-1997	37.069	-76.55	1	1.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0982	25-AUG-1997	37.053	-76.556	1	9.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0983	25-AUG-1997	37.044	-76.548	1	8.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0984	25-AUG-1997	36.993	-76.472	1	8.4	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0985	25-AUG-1997	37.004	-76.329	1	2.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0986	25-AUG-1997	36.992	-76.515	1	2.3	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0987	25-AUG-1997	36.979	-76.447	1	9.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0988	25-AUG-1997	36.975	-76.369	1	3.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0989	25-AUG-1997	36.954	-76.278	1	3.0	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0990	25-AUG-1997	36.917	-76.413	1	2.7	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0991	25-AUG-1997	36.912	-76.413	1	2.6	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0992	25-AUG-1997	36.895	-76.466	1	4.8	m	
EMAP Mid-Atlantic Integrated Assessment/Chesapeake Bay Program	1997	MA97-0993	25-AUG-1997	36.885	-76.456	1	1.2	m	
EMAP Mid-Atlantic Integrated Assessment/National Park Service	1998	MA98-0002	08-OCT-1998	38.247	-75.149	1	2.8	m	
EMAP Mid-Atlantic Integrated Assessment/National Park Service	1998	MA98-0003	06-OCT-1998	38.239	-75.209	1	1.3	m	
EMAP Mid-Atlantic Integrated Assessment/National Park Service	1998	MA98-0006	07-OCT-1998	38.107	-75.235	1	1.9	m	
EMAP Mid-Atlantic Integrated Assessment/National Park Service	1998	MA98-0009	06-OCT-1998	38.004	-75.386	1	1.7	m	
EMAP Mid-Atlantic Integrated Assessment/National Park Service	1998	MA98-0014	07-OCT-1998	38.067	-75.331	1	1.5	m	
EMAP Mid-Atlantic Integrated Assessment/National Park Service	1998	MA98-0018	05-OCT-1998	38.285	-75.131	1	1.9	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0032	15-AUG-1998	38.228	-75.175	1	1.5	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0046	12-AUG-1998	37.375	-75.754	1	7.8	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0050	15-AUG-1998	37.884	-75.394	1	0.9	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0055	11-AUG-1998	37.211	-75.92	1	1.3	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0056	11-AUG-1998	37.333	-75.892	1	4.3	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0058	13-AUG-1998	37.458	-75.678	1	10.4	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0067	01-AUG-1998	37.336	-76.4	1	2.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0073	22-AUG-1998	38.567	-76.207	1	2.3	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0074	24-AUG-1998	38.745	-76.25	1	4.2	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0078	30-AUG-1998	38.929	-76.315	1	2.2	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0079	13-JUL-1998	39.507	-75.915	1	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0080	01-AUG-1998	37.483	-76.275	1	0.8	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0081	14-AUG-1998	37.848	-75.686	1	2.8	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0083	10-AUG-1998	37.419	-75.961	1	1.3	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0086	20-AUG-1998	38.115	-75.888	1	1.6	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0088	13-AUG-1998	37.552	-75.889	1	2.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0089	15-JUL-1998	39.214	-76.452	1	2.3	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0090	15-JUL-1998	39.249	-76.553	1	9.9	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0091	30-JUL-1998	37.522	-76.412	1	8.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0093	27-JUL-1998	38.132	-76.482	1	2.7	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0097	30-AUG-1998	38.877	-76.126	1	4.3	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0118	16-JUL-1998	39.047	-76.555	1	7.5	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0144	16-JUL-1998	38.951	-76.538	1	5.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0171	04-AUG-1998	37.566	-76.883	1	2.9	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0231	10-AUG-1998	37.28	-76.008	1	1.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0253	19-AUG-1998	38.043	-75.662	1	4.4	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0313	13-JUL-1998	39.527	-76.07	1	1.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0322	31-AUG-1998	39.36	-76.145	1	8.4	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0356	17-SEP-1998	39.045	-76.396	1	8.4	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0376	23-AUG-1998	38.701	-75.991	1	2.2	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0378	18-JUL-1998	38.675	-77.113	1	1.5	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0381	14-SEP-1998	38.648	-76.497	1	10.2	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0383	23-AUG-1998	38.604	-76.113	1	4.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0391	22-AUG-1998	38.534	-76.325	1	3.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0392	20-JUL-1998	38.506	-76.668	1	2.8	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0394	23-JUL-1998	38.467	-77.296	1	3.2	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0437	05-SEP-1998	39.583	-75.49	1	2.7	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0440	05-SEP-1998	39.571	-75.535	1	2.4	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0447	04-SEP-1998	39.447	-75.506	1	2.4	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0451	03-SEP-1998	39.383	-75.333	1	4.6	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0452	04-SEP-1998	39.381	-75.435	1	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0454	04-SEP-1998	39.346	-75.481	1	2.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0457	02-SEP-1998	39.24	-75.424	1	6.5	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0460	19-SEP-1998	39.178	-75.353	1	4.3	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0465	19-SEP-1998	39.129	-75.251	1	5.1	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0843	22-JUL-1998	38.391	-76.521	1	7.4	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0846	24-JUL-1998	38.356	-77.22	1	5.9	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0859	22-JUL-1998	38.298	-76.435	1	9.2	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0864	25-JUL-1998	38.219	-76.846	1	7.1	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0872	21-AUG-1998	38.168	-76.001	1	3.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0873	28-JUL-1998	38.148	-77.083	1	4.5	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0874	13-SEP-1998	38.151	-76.121	1	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0877	25-JUL-1998	38.102	-76.57	1	7.2	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0881	20-AUG-1998	38.065	-75.896	1	7.5	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0899	13-SEP-1998	37.915	-76.151	1	26.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0915	29-JUL-1998	37.694	-76.573	1	5.1	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0918	12-SEP-1998	37.681	-75.927	1	5.8	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0926	30-JUL-1998	37.611	-76.41	1	9.2	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0928	12-SEP-1998	37.591	-76.049	1	14.2	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0932	12-SEP-1998	37.52	-76.271	1	4.8	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0944	11-SEP-1998	37.378	-76.026	1	11.5	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0945	03-AUG-1998	37.369	-76.645	1	3.5	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0951	08-AUG-1998	37.316	-77.223	1	9.3	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0959	10-SEP-1998	37.276	-76.322	1	4.7	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0961	03-AUG-1998	37.249	-76.523	1	10.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0966	07-AUG-1998	37.23	-76.809	1	2.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0971	07-AUG-1998	37.212	-76.901	1	7.2	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0973	06-AUG-1998	37.184	-76.738	1	7.6	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0976	11-SEP-1998	37.143	-76.196	1	11.2	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0985	05-AUG-1998	37.003	-76.329	1	3.2	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-0988	05-AUG-1998	36.975	-76.369	1	4.8	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-1021	27-AUG-1998	38.934	-76.223	1	3.5	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-1022	29-AUG-1998	38.868	-76.271	1	12.3	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-1023	27-AUG-1998	38.898	-76.24	1	1.4	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-1024	29-AUG-1998	38.851	-76.349	1	3.7	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-1025	29-AUG-1998	38.871	-76.303	1	5.6	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-1026	27-AUG-1998	38.85	-76.212	1	3.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-1027	26-AUG-1998	38.825	-76.246	1	1.6	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-1028	26-AUG-1998	38.834	-76.235	1	12.3	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-1029	26-AUG-1998	38.799	-76.196	1	2.9	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-1030	26-AUG-1998	38.797	-76.204	1	6.6	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-1061	31-AUG-1998	39.005	-76.254	1	6.0	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-1064	18-SEP-1998	39.266	-75.323	1	6.4	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-1066	28-JUL-1998	37.99	-76.902	1	3.3	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-1067	27-JUL-1998	38.065	-76.375	1	4.6	m	
EMAP Mid-Atlantic Integrated Assessment/USEPA Office of Research and Development	1998	MA98-1068	06-AUG-1998	37.073	-76.574	1	2.8	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0001	15-AUG-2000	38.238	-75.207	1	1.7	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0002	15-AUG-2000	38.256	-75.192	1	1.4	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0003	15-AUG-2000	38.146	-75.284	1	1.2	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0004	15-AUG-2000	38.066	-75.33	1	1.8	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0005	15-AUG-2000	38.074	-75.359	1	1.4	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0006	15-AUG-2000	38.036	-75.268	1	2.2	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0007	15-AUG-2000	38.108	-75.229	1	1.9	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0008	16-AUG-2000	38.215	-75.178	1	2.0	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0009	16-AUG-2000	38.246	-75.149	1	2.4	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0010	16-AUG-2000	38.294	-75.124	1			
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0011	16-AUG-2000	38.32	-75.107	1			
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0012	16-AUG-2000	38.327	-75.104	1	2.1	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0013	24-AUG-2000	38.193	-75.232	1	1.9	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0014	24-AUG-2000	38.222	-75.221	1	1.7	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0015	24-AUG-2000	38.246	-75.203	1	1.6	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0022	24-AUG-2000	38.295	-75.162	1	1.3	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0024	24-AUG-2000	38.268	-75.199	1	1.0	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0025	24-AUG-2000	38.286	-75.207	1	1.2	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0027	17-AUG-2000	38.392	-75.12	1	2.0	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0028	17-AUG-2000	38.395	-75.129	1	1.5	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0029	17-AUG-2000	38.404	-75.147	1	1.5	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0030	17-AUG-2000	38.411	-75.171	1	1.1	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0031	17-AUG-2000	38.424	-75.189	1	1.0	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0032	17-AUG-2000	38.414	-75.185	1	1.1	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0033	17-AUG-2000	38.408	-75.175	1	1.2	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0034	17-AUG-2000	38.408	-75.186	1	1.1	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0038	17-AUG-2000	38.355	-75.147	1	0.6	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0039	17-AUG-2000	38.357	-75.168	1			
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0040	17-AUG-2000	38.34	-75.13	1	1.4	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0041	15-AUG-2000	38.334	-75.09	1			
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0042	14-AUG-2000	38.355	-75.089	1			
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0043	14-AUG-2000	38.373	-75.103	1			
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0044	16-AUG-2000	38.389	-75.092	1			
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0045	16-AUG-2000	38.413	-75.09	1			
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0046	16-AUG-2000	38.428	-75.105	1			
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0047	16-AUG-2000	38.442	-75.078	1			
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0048	15-AUG-2000	38.359	-75.131	1			
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0049	15-AUG-2000	38.373	-75.135	1			
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0050	17-AUG-2000	38.454	-75.138	1			
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0051	16-AUG-2000	38.458	-75.09	1			
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0052	16-AUG-2000	38.453	-75.064	1			
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0053	03-AUG-2000	38.168	-75.237	1			
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0054	02-AUG-2000	38.099	-75.275	1			
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0055	02-AUG-2000	38.135	-75.251	1			
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2000	MD00-0056	01-AUG-2000	38.022	-75.333	1			
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0001	15-AUG-2001	38.238	-75.207	2	1.4	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0002	15-AUG-2001	38.256	-75.192	2	1.1	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0003	15-AUG-2001	38.146	-75.284	2	0.8	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0004	15-AUG-2001	38.066	-75.33	2	1.5	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0005	15-AUG-2001	38.074	-75.359	2	1.1	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0006	15-AUG-2001	38.036	-75.268	2	1.9	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0007	15-AUG-2001	38.108	-75.229	2	1.5	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0008	16-AUG-2001	38.215	-75.178	2	2.0	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0009	16-AUG-2001	38.246	-75.149	2	2.1	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0010	16-AUG-2001	38.294	-75.124	2	1.7	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0011	16-AUG-2001	38.32	-75.107	2	2.3	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0012	16-AUG-2001	38.327	-75.104	2	1.1	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0013	23-AUG-2001	38.193	-75.232	2	2.0	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0014	23-AUG-2001	38.222	-75.221	2	1.7	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0015	23-AUG-2001	38.246	-75.203	2	1.6	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0016	23-AUG-2001	38.296	-75.18	2	0.6	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0022	23-AUG-2001	38.295	-75.162	2	1.8	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0024	23-AUG-2001	38.268	-75.199	2	1.0	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0025	23-AUG-2001	38.286	-75.207	2	0.9	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0027	22-AUG-2001	38.392	-75.12	2	1.8	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0028	22-AUG-2001	38.395	-75.129	2	1.5	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0029	22-AUG-2001	38.404	-75.147	2	1.2	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0030	22-AUG-2001	38.411	-75.171	2	1.0	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0031	22-AUG-2001	38.424	-75.189	2	0.9	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0032	22-AUG-2001	38.414	-75.185	2	1.0	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0033	22-AUG-2001	38.408	-75.175	2	1.1	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0034	22-AUG-2001	38.408	-75.186	2	0.9	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0038	22-AUG-2001	38.355	-75.147	2	0.5	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0039	22-AUG-2001	38.357	-75.168	2			
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0040	22-AUG-2001	38.34	-75.13	2	1.7	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0041	09-AUG-2001	38.334	-75.09	2	7.5	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0042	09-AUG-2001	38.355	-75.089	2	4.2	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0043	09-AUG-2001	38.373	-75.103	2	2.0	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0044	09-AUG-2001	38.389	-75.092	2	2.4	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0045	09-AUG-2001	38.413	-75.09	2	2.1	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0046	09-AUG-2001	38.428	-75.105	2	1.5	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0047	09-AUG-2001	38.442	-75.078	2	1.8	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0048	09-AUG-2001	38.359	-75.131	2	1.3	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0049	09-AUG-2001	38.373	-75.135	2	6.4	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0050	09-AUG-2001	38.454	-75.138	2			
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0051	09-AUG-2001	38.458	-75.09	2	1.1	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0052	09-AUG-2001	38.453	-75.064	2			
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0053	23-AUG-2001	38.168	-75.237	2	1.8	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0054	23-AUG-2001	38.099	-75.275	2	1.8	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0055	23-AUG-2001	38.135	-75.251	2	1.7	m	
National Coastal Assessment-Southeast/Maryland Dept. of Natural Resouces-Coastal Bays	2001	MD01-0056	23-AUG-2001	38.022	-75.333	2	1.8	m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0001-A	03-AUG-2005	38.082	-75.22	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0001-A	25-AUG-2005	38.082	-75.22	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0002-A	21-SEP-2005	38.639	-76.199	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0003-B	19-SEP-2005	38.305	-76.964	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0003-B	30-SEP-2005	38.305	-76.964	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0004-A	04-AUG-2005	38.169	-75.233	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0004-A	25-AUG-2005	38.169	-75.233	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0005-A	30-AUG-2005	38.2	-76.255	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0005-A	12-SEP-2005	38.2	-76.255	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0007-A	24-AUG-2005	38.35	-75.091	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0008-A	08-SEP-2005	39.005	-76.504	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0009-B	14-SEP-2005	38.217	-75.85	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0009-B	20-SEP-2005	38.217	-75.85	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0010-A	30-AUG-2005	38.26	-76.279	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0010-A	12-SEP-2005	38.26	-76.279	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0011-A	19-SEP-2005	38.336	-76.84	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0011-A	29-SEP-2005	38.336	-76.84	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0012-A	03-AUG-2005	38.078	-75.349	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0012-A	25-AUG-2005	38.078	-75.349	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0013-A	30-AUG-2005	38.026	-76.137	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0013-A	09-SEP-2005	38.026	-76.137	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0014-A	28-SEP-2005	38.913	-76.291	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0015-B	01-SEP-2005	39.437	-76.059	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0016-A	21-SEP-2005	38.888	-76.111	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0017-A	30-AUG-2005	38.088	-76.208	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0017-A	12-SEP-2005	38.088	-76.208	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0018-B	31-AUG-2005	39.209	-76.522	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0018-B	11-SEP-2005	39.209	-76.522	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0019-A	14-SEP-2005	38.111	-75.875	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0019-A	28-SEP-2005	38.111	-75.875	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0020-A	10-SEP-2005	38.838	-76.478	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0020-A	13-SEP-2005	38.838	-76.478	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0021-A	29-AUG-2005	38.236	-76.35	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0021-A	12-SEP-2005	38.236	-76.35	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0022-A	04-AUG-2005	38.187	-75.204	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0022-A	24-AUG-2005	38.187	-75.204	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0023-A	10-SEP-2005	38.505	-76.483	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0023-A	13-SEP-2005	38.505	-76.483	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0024-A	03-AUG-2005	38.101	-75.322	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0024-A	25-AUG-2005	38.101	-75.322	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0025-A	29-AUG-2005	38.101	-76.494	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2005	MD05-0025-A	12-SEP-2005	38.101	-76.494	1		m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2006	MD06-0026-A	26-SEP-2006	38.243	-76.801	1	2.7	m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2006	MD06-0027-A	08-SEP-2006	39.124	-76.42	1	4.0	m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2006	MD06-0028-A	06-SEP-2006	37.96	-76.085	1	6.0	m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2006	MD06-0028-A	22-SEP-2006	37.96	-76.085	2	6.0	m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2006	MD06-0029-A	07-SEP-2006	38.659	-76.391	1	12.0	m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2006	MD06-0029-A	22-SEP-2006	38.659	-76.391	2	12.0	m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2006	MD06-0030-A	09-SEP-2006	38.048	-76.436	1	13.0	m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2006	MD06-0030-A	21-SEP-2006	38.048	-76.436	2	13.0	m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2006	MD06-0031-A	07-SEP-2006	38.41	-76.391	1	12.5	m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2006	MD06-0031-A	20-SEP-2006	38.41	-76.391	2	12.5	m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2006	MD06-0032-A	07-SEP-2006	38.582	-76.452	1	12.0	m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2006	MD06-0032-A	20-SEP-2006	38.582	-76.452	2	12.0	m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2006	MD06-0033-A	02-AUG-2006	38.043	-75.283	1	1.5	m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2006	MD06-0034-A	09-SEP-2006	37.978	-76.402	1	6.0	m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2006	MD06-0034-A	21-SEP-2006	37.978	-76.402	2	6.0	m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2006	MD06-0035-C	08-SEP-2006	39.262	-76.304	1	4.4	m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2006	MD06-0036-A	01-AUG-2006	38.44	-75.088	1	0.5	m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2006	MD06-0037-A	12-SEP-2006	39.03	-76.199	1	5.1	m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2006	MD06-0038-A	11-SEP-2006	38.451	-77.288	1	5.1	m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2006	MD06-0039-A	02-AUG-2006	38.197	-75.246	1	1.0	m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2006	MD06-0040-A	07-SEP-2006	38.592	-76.415	1	15.0	m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2006	MD06-0040-A	22-SEP-2006	38.592	-76.415	2	15.0	m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2006	MD06-0041-A	02-AUG-2006	38.142	-75.231	1	2.0	m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2006	MD06-0042-B	14-SEP-2006	38.665	-75.953	1	2.7	m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2006	MD06-0043-A	07-SEP-2006	38.443	-76.323	1	3.0	m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2006	MD06-0043-A	22-SEP-2006	38.443	-76.323	2	3.0	m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2006	MD06-0044-A	21-SEP-2006	38.283	-76.952	1	10.0	m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2006	MD06-0045-A	01-AUG-2006	38.361	-75.104	1	1.5	m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2006	MD06-0046-B	22-SEP-2006	38.267	-76.123	1	3.0	m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2006	MD06-0047-A	06-SEP-2006	38.961	-76.47	1	1.6	m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2006	MD06-0047-A	07-SEP-2006	38.961	-76.47	2	1.6	m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2006	MD06-0048-A	07-SEP-2006	39.441	-75.979	2	1.6	m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2006	MD06-0049-A	28-SEP-2006	38.865	-76.199	1	1.5	m	
National Coastal Assessment-Northeast/Chesapeake Bay Program	2006	MD06-0050-A	22-SEP-2006	38.227	-76.011	1	3.0	m	
R-EMAP Region 2 1993-94	1993	NB018	10-AUG-1993	40.727	-74.101	1	9.4	m	
R-EMAP Region 2 1993-94	1993	NB021	26-AUG-1993	40.712	-74.12	1	2.1	m	
R-EMAP Region 2 1993-94	1993	NB025	11-AUG-1993	40.704	-74.116	1	4.3	m	
R-EMAP Region 2 1993-94	1993	NB027	11-AUG-1993	40.698	-74.122	1	4.3	m	
R-EMAP Region 2 1993-94	1993	NB036	26-AUG-1993	40.675	-74.128	1	2.8	m	
R-EMAP Region 2 1993-94	1993	NB039	13-AUG-1993	40.674	-74.128	1	3.4	m	
R-EMAP Region 2 1993-94	1993	NB044	13-AUG-1993	40.655	-74.156	1	3.5	m	
R-EMAP Region 2 1993-94	1993	NB045	04-AUG-1993	40.65	-74.146	1	12.8	m	
R-EMAP Region 2 1993-94	1993	NB047	03-AUG-1993	40.64	-74.192	1	11.3	m	
R-EMAP Region 2 1993-94	1993	NB052	04-AUG-1993	40.647	-74.154	1	14.0	m	
R-EMAP Region 2 1993-94	1993	NB053	05-AUG-1993	40.645	-74.149	1	14.0	m	
R-EMAP Region 2 1993-94	1993	NB065	26-AUG-1993	40.717	-74.108	1	4.0	m	
R-EMAP Region 2 1993-94	1993	NB066	11-AUG-1993	40.718	-74.122	1	6.1	m	
R-EMAP Region 2 1993-94	1993	NB075	13-AUG-1993	40.528	-74.25	1	5.5	m	
R-EMAP Region 2 1993-94	1994	NB102	18-AUG-1994	40.688	-74.158	1	12.8	m	
R-EMAP Region 2 1993-94	1994	NB103	05-AUG-1994	40.662	-74.136	1	3.4	m	
R-EMAP Region 2 1993-94	1994	NB104	05-AUG-1994	40.712	-74.111	1	4.6	m	
R-EMAP Region 2 1993-94	1994	NB105	18-AUG-1994	40.686	-74.129	1	13.1	m	
R-EMAP Region 2 1993-94	1994	NB106	25-AUG-1994	40.667	-74.13	1	3.4	m	
R-EMAP Region 2 1993-94	1994	NB107	16-SEP-1994	40.555	-74.237	1	4.6	m	
R-EMAP Region 2 1993-94	1994	NB108	23-AUG-1994	40.74	-74.118	1	7.3	m	
R-EMAP Region 2 1993-94	1994	NB109	21-SEP-1994	40.614	-74.197	1	2.1	m	
R-EMAP Region 2 1993-94	1994	NB110	19-SEP-1994	40.696	-74.115	1	3.7	m	
R-EMAP Region 2 1993-94	1994	NB111	24-AUG-1994	40.721	-74.121	1	4.3	m	
R-EMAP Region 2 1993-94	1994	NB112	24-AUG-1994	40.681	-74.141	1	13.1	m	
R-EMAP Region 2 1993-94	1994	NB113	20-SEP-1994	40.651	-74.157	1	3.0	m	
R-EMAP Region 2 1993-94	1994	NB114	23-AUG-1994	40.736	-74.16	1	6.1	m	
R-EMAP Region 2 1993-94	1994	NB115	19-SEP-1994	40.649	-74.106	1	12.5	m	
R-EMAP Region 2 1998	1998	NB201	01-JUL-1998	40.665	-74.141	1			
R-EMAP Region 2 1998	1998	NB201	15-AUG-1998	40.665	-74.141	2	13.4	m	
R-EMAP Region 2 1998	1998	NB202	01-JUL-1998	40.646	-74.177	1			
R-EMAP Region 2 1998	1998	NB202	17-AUG-1998	40.646	-74.177	2	11.3	m	
R-EMAP Region 2 1998	1998	NB203	01-JUL-1998	40.615	-74.202	1			
R-EMAP Region 2 1998	1998	NB203	16-JUL-1998	40.615	-74.202	2	2.1	m	
R-EMAP Region 2 1998	1998	NB204	01-JUL-1998	40.615	-74.202	1			
R-EMAP Region 2 1998	1998	NB204	16-JUL-1998	40.615	-74.202	2	13.4	m	
R-EMAP Region 2 1998	1998	NB205	20-AUG-1998	40.738	-74.117	1	6.7	m	
R-EMAP Region 2 1998	1999	NB205	01-JUL-1999	40.738	-74.117	2			
R-EMAP Region 2 1998	1998	NB206	18-AUG-1998	40.677	-74.139	1	12.5	m	
R-EMAP Region 2 1998	1999	NB206	01-JUL-1999	40.677	-74.139	2			
R-EMAP Region 2 1998	1998	NB207	13-JUL-1998	40.648	-74.115	1	7.0	m	
R-EMAP Region 2 1998	1999	NB207	01-JUL-1999	40.648	-74.115	2			
R-EMAP Region 2 1998	1998	NB208	13-AUG-1998	40.535	-74.252	1	11.3	m	
R-EMAP Region 2 1998	1999	NB208	01-JUL-1999	40.535	-74.252	2			
R-EMAP Region 2 1998	1998	NB209	14-AUG-1998	40.553	-74.245	1	11.9	m	
R-EMAP Region 2 1998	1999	NB209	01-JUL-1999	40.553	-74.245	2			
R-EMAP Region 2 1998	1998	NB210	18-JUL-1998	40.559	-74.216	1	11.9	m	
R-EMAP Region 2 1998	1999	NB210	01-JUL-1999	40.559	-74.216	2			
R-EMAP Region 2 1998	1998	NB211	17-AUG-1998	40.638	-74.194	1	11.3	m	
R-EMAP Region 2 1998	1999	NB211	01-JUL-1999	40.638	-74.194	2			
R-EMAP Region 2 1998	1998	NB212	15-AUG-1998	40.669	-74.138	1	14.0	m	
R-EMAP Region 2 1998	1999	NB212	01-JUL-1999	40.669	-74.138	2			
R-EMAP Region 2 1998	1998	NB213	15-AUG-1998	40.644	-74.164	1	5.5	m	
R-EMAP Region 2 1998	1999	NB213	01-JUL-1999	40.664	-74.164	2			
R-EMAP Region 2 1998	1998	NB214	18-JUL-1998	40.58	-74.208	1	4.9	m	
R-EMAP Region 2 1998	1999	NB214	01-JUL-1999	40.58	-74.208	2			
R-EMAP Region 2 1998	1998	NB216	17-AUG-1998	40.688	-74.136	1	13.7	m	
R-EMAP Region 2 1998	1999	NB216	01-JUL-1999	40.688	-74.136	2			
R-EMAP Region 2 1998	1998	NB217	11-JUL-1998	40.692	-74.119	1	4.0	m	
R-EMAP Region 2 1998	1999	NB217	01-JUL-1999	40.692	-74.119	2			
R-EMAP Region 2 1998	1998	NB218	16-JUL-1998	40.645	-74.127	1	9.8	m	
R-EMAP Region 2 1998	1999	NB218	01-JUL-1999	40.645	-74.127	2			
R-EMAP Region 2 1998	1998	NB219	18-JUL-1998	40.559	-74.233	1	9.4	m	
R-EMAP Region 2 1998	1999	NB219	01-JUL-1999	40.559	-74.233	2			
R-EMAP Region 2 1998	1998	NB222	11-JUL-1998	40.654	-74.142	1	3.0	m	
R-EMAP Region 2 1998	1999	NB222	01-JUL-1999	40.654	-74.142	2			
R-EMAP Region 2 1998	1998	NB223	15-AUG-1998	40.65	-74.166	1	3.0	m	
R-EMAP Region 2 1998	1999	NB223	01-JUL-1999	40.65	-74.166	2			
R-EMAP Region 2 1998	1998	NB224	16-JUL-1998	40.606	-74.203	1	13.1	m	
R-EMAP Region 2 1998	1999	NB224	01-JUL-1999	40.606	-74.203	2			
R-EMAP Region 2 1998	1998	NB225	20-AUG-1998	40.724	-74.101	1	10.4	m	
R-EMAP Region 2 1998	1999	NB225	01-JUL-1999	40.724	-74.101	2			
R-EMAP Region 2 1998	1998	NB226	11-JUL-1998	40.673	-74.131	1	2.7	m	
R-EMAP Region 2 1998	1999	NB226	01-JUL-1999	40.673	-74.131	2			
R-EMAP Region 2 1998	1998	NB227	18-AUG-1998	40.704	-74.117	1	11.9	m	
R-EMAP Region 2 1998	1999	NB227	01-JUL-1999	40.704	-74.117	2			
R-EMAP Region 2 1998	1998	NB228	13-JUL-1998	40.646	-74.102	1	14.3	m	
R-EMAP Region 2 1998	1999	NB228	01-JUL-1999	40.646	-74.102	2			
R-EMAP Region 2 1998	1998	NB229	14-AUG-1998	40.516	-74.255	1	10.1	m	
R-EMAP Region 2 1998	1999	NB229	01-JUL-1999	40.516	-74.255	2			
R-EMAP Region 2 1998	1998	NB230	21-AUG-1998	40.545	-74.249	1	5.5	m	
R-EMAP Region 2 1998	1999	NB230	01-JUL-1999	40.545	-74.249	2			
R-EMAP Region 2 1998	1998	NB231	21-AUG-1998	40.66	-74.138	1	3.4	m	
R-EMAP Region 2 1998	1999	NB231	01-JUL-1999	40.66	-74.138	2			
R-EMAP Region 2 2003	2003	NB301	26-AUG-2003	40.66	-74.138	1	14.3	m	
R-EMAP Region 2 2003	2003	NB301	27-AUG-2003	40.66	-74.138	2	14.3	m	
R-EMAP Region 2 2003	2003	NB305	30-AUG-2003	40.665	-74.141	1	8.4	m	
R-EMAP Region 2 2003	2003	NB305	02-SEP-2003	40.665	-74.141	2	8.4	m	
R-EMAP Region 2 2003	2003	NB306	15-JUL-2003	40.669	-74.138	1	8.5	m	
R-EMAP Region 2 2003	2003	NB306	16-JUL-2003	40.669	-74.138	2	8.5	m	
R-EMAP Region 2 2003	2003	NB307	16-JUL-2003	40.643	-74.143	1	5.8	m	
R-EMAP Region 2 2003	2003	NB307	17-JUL-2003	40.643	-74.143	2	5.8	m	
R-EMAP Region 2 2003	2003	NB309	04-SEP-2003	40.644	-74.164	1	10.4	m	
R-EMAP Region 2 2003	2003	NB309	05-SEP-2003	40.644	-74.164	2	10.4	m	
R-EMAP Region 2 2003	2003	NB310	17-JUL-2003	40.649	-74.167	1	11.3	m	
R-EMAP Region 2 2003	2003	NB310	18-JUL-2003	40.649	-74.167	2	11.3	m	
R-EMAP Region 2 2003	2003	NB312	26-AUG-2003	40.649	-74.159	1	14.6	m	
R-EMAP Region 2 2003	2003	NB312	27-AUG-2003	40.649	-74.159	2	14.6	m	
R-EMAP Region 2 2003	2003	NB313	10-SEP-2003	40.614	-74.201	1	2.7	m	
R-EMAP Region 2 2003	2003	NB313	12-SEP-2003	40.614	-74.201	2	2.7	m	
R-EMAP Region 2 2003	2003	NB314	16-JUL-2003	40.581	-74.208	1	4.3	m	
R-EMAP Region 2 2003	2003	NB314	17-JUL-2003	40.581	-74.208	2	4.3	m	
R-EMAP Region 2 2003	2003	NB316	27-AUG-2003	40.606	-74.205	1	12.8	m	
R-EMAP Region 2 2003	2003	NB318	05-SEP-2003	40.591	-74.203	1	11.6	m	
R-EMAP Region 2 2003	2003	NB318	09-SEP-2003	40.591	-74.203	2	11.6	m	
R-EMAP Region 2 2003	2003	NB319	04-SEP-2003	40.724	-74.101	1	9.5	m	
R-EMAP Region 2 2003	2003	NB319	05-SEP-2003	40.724	-74.101	2	9.5	m	
R-EMAP Region 2 2003	2003	NB323	04-SEP-2003	40.718	-74.123	1	2.4	m	
R-EMAP Region 2 2003	2003	NB323	05-SEP-2003	40.718	-74.123	2	2.4	m	
R-EMAP Region 2 2003	2003	NB324	16-JUL-2003	40.738	-74.117	1	10.7	m	
R-EMAP Region 2 2003	2003	NB324	17-JUL-2003	40.738	-74.117	2	10.7	m	
R-EMAP Region 2 2003	2003	NB325	30-AUG-2003	40.688	-74.135	1	11.0	m	
R-EMAP Region 2 2003	2003	NB325	02-SEP-2003	40.688	-74.135	2	11.0	m	
R-EMAP Region 2 2003	2003	NB326	15-JUL-2003	40.674	-74.131	1	2.9	m	
R-EMAP Region 2 2003	2003	NB326	16-JUL-2003	40.674	-74.131	2	2.9	m	
R-EMAP Region 2 2003	2003	NB327	30-AUG-2003	40.677	-74.138	1	11.0	m	
R-EMAP Region 2 2003	2003	NB327	02-SEP-2003	40.677	-74.138	2	11.0	m	
R-EMAP Region 2 2003	2003	NB329	18-JUL-2003	40.705	-74.117	1	10.7	m	
R-EMAP Region 2 2003	2003	NB329	18-AUG-2003	40.705	-74.117	2	10.7	m	
R-EMAP Region 2 2003	2003	NB330	03-SEP-2003	40.749	-74.082	1	4.9	m	
R-EMAP Region 2 2003	2003	NB330	04-SEP-2003	40.749	-74.082	2	4.9	m	
R-EMAP Region 2 2003	2003	NB330	05-SEP-2003	40.749	-74.082	3	4.9	m	
R-EMAP Region 2 2003	2003	NB331	15-JUL-2003	40.648	-74.115	1	2.9	m	
R-EMAP Region 2 2003	2003	NB331	16-JUL-2003	40.648	-74.115	2	2.9	m	
R-EMAP Region 2 2003	2003	NB350	10-SEP-2003	40.645	-74.126	1	4.0	m	
R-EMAP Region 2 2003	2003	NB350	12-SEP-2003	40.645	-74.126	2	4.0	m	
R-EMAP Region 2 2003	2003	NB352	26-AUG-2003	40.648	-74.092	1	2.4	m	
R-EMAP Region 2 2003	2003	NB352	27-AUG-2003	40.648	-74.092	2	2.4	m	
R-EMAP Region 2 2003	2003	NB353	02-SEP-2003	40.559	-74.234	1	13.7	m	
R-EMAP Region 2 2003	2003	NB353	04-SEP-2003	40.559	-74.234	2	13.7	m	
R-EMAP Region 2 2003	2003	NB354	30-AUG-2003	40.517	-74.256	1	3.4	m	
R-EMAP Region 2 2003	2003	NB354	02-SEP-2003	40.517	-74.256	2	3.4	m	
R-EMAP Region 2 2003	2003	NB355	17-JUL-2003	40.553	-74.247	1	1.7	m	
R-EMAP Region 2 2003	2003	NB355	18-JUL-2003	40.553	-74.247	2	1.7	m	
R-EMAP Region 2 2003	2003	NB357	02-SEP-2003	40.532	-74.245	1	9.5	m	
R-EMAP Region 2 2003	2003	NB357	04-SEP-2003	40.532	-74.245	2	9.5	m	
R-EMAP Region 2 2003	2003	NB359	03-SEP-2003	40.545	-74.249	1	5.5	m	
R-EMAP Region 2 2003	2003	NB359	04-SEP-2003	40.545	-74.249	2	5.5	m	
R-EMAP Region 2 2003	2003	NB360	05-SEP-2003	40.559	-74.217	1	2.7	m	
R-EMAP Region 2 2003	2003	NB360	09-SEP-2003	40.559	-74.217	2	2.7	m	
R-EMAP Region 2 2003	2003	NB361	03-SEP-2003	40.74	-74.141	1	11.6	m	
R-EMAP Region 2 2003	2003	NB361	04-SEP-2003	40.74	-74.141	2	11.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0001-A	22-AUG-2000	40.485	-74.341	1	14.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0003-B	15-AUG-2000	40.435	-74.038	1	4.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0005-A	22-AUG-2000	40.506	-74.314	1	8.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0007-A	10-AUG-2000	40.476	-74.071	1	7.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0009-A	10-AUG-2000	40.661	-74.14	1	10.4	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0011-B	21-AUG-2000	40.762	-74.161	1	5.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0013-A	21-AUG-2000	40.805	-74.14	1	5.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0015-A	16-AUG-2000	40.923	-73.919	1	10.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0017-A	12-SEP-2000	38.992	-74.833	1	0.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0019-A	31-AUG-2000	39.091	-74.739	1	6.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0021-A	31-AUG-2000	39.121	-74.718	1	6.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0023-A	31-AUG-2000	39.204	-74.655	1	3.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0025-A	12-SEP-2000	39.292	-74.62	1	9.4	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0027-A	11-SEP-2000	39.365	-74.716	1	2.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0029-A	08-SEP-2000	39.37	-74.477	1	2.1	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0031-A	11-SEP-2000	39.449	-74.724	1	1.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0033-A	08-SEP-2000	39.444	-74.454	1	0.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0035-A	07-SEP-2000	39.505	-74.399	1	2.1	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0037-A	07-SEP-2000	39.594	-74.551	1	2.1	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0039-A	06-SEP-2000	39.554	-74.315	1	1.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0041-A	07-SEP-2000	39.612	-74.589	1	4.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0043-A	06-SEP-2000	39.64	-74.205	1	2.1	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0045-A	05-SEP-2000	39.743	-74.148	1	2.8	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0047-A	05-SEP-2000	39.81	-74.102	1	1.1	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0049-A	29-AUG-2000	39.933	-74.141	1	2.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0051-A	29-AUG-2000	39.99	-74.074	1	1.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0053-A	28-AUG-2000	40.092	-74.078	1	1.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0055-A	28-AUG-2000	40.187	-74.02	1	4.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0057-A	22-AUG-2000	40.348	-74.081	1	1.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0059-A	15-AUG-2000	40.378	-74.024	1	3.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0061-A	03-OCT-2000	38.972	-74.982	1	7.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0063-A	12-OCT-2000	39.13	-75.121	1	4.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0065-A	12-OCT-2000	39.201	-75.221	1	5.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0067-A	03-OCT-2000	39.163	-74.9	1	1.1	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0069-A	12-OCT-2000	39.248	-75.208	1	3.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0071-A	13-OCT-2000	39.32	-75.334	1	5.5	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0073-A	10-OCT-2000	40.079	-74.87	1	13.4	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0075-A	10-OCT-2000	39.983	-75.067	1	13.4	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0077-A	10-OCT-2000	39.88	-75.179	1	10.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0079-A	11-OCT-2000	39.845	-75.338	1	12.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0081-A	04-OCT-2000	39.083	-75.183	1	14.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0083-B	13-SEP-2000	38.967	-74.952	1	1.5	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0085-A	13-SEP-2000	38.963	-74.926	1	2.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0087-A	14-SEP-2000	39.174	-74.859	1	5.1	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0089-A	15-SEP-2000	39.204	-75.031	1	2.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0091-A	20-SEP-2000	39.346	-75.358	1	2.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0093-A	15-SEP-2000	39.347	-75.024	1	2.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0095-C	19-SEP-2000	39.502	-75.508	1	1.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0097-A	20-SEP-2000	39.392	-75.227	1	5.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	NJ00-0101-B	21-SEP-2000	39.626	-75.449	1	0.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0002-A	30-AUG-2001	40.472	-74.097	1	6.8	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0006-A	25-SEP-2001	40.482	-74.24	1	4.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0008-A	29-AUG-2001	40.522	-73.97	1	4.8	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0010-C	29-AUG-2001	40.684	-74.041	1	13.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0012-A	29-OCT-2001	40.706	-74.108	1	0.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0014-B	28-AUG-2001	40.842	-73.959	1	8.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0016-A	12-SEP-2001	38.95	-74.903	1	2.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0018-A	12-SEP-2001	39.01	-74.842	1	1.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0020-A	30-AUG-2001	39.095	-74.785	1	1.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0022-A	30-AUG-2001	39.187	-74.671	1	4.4	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0024-A	27-SEP-2001	39.296	-74.753	1	2.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0026-A	18-JUL-2001	39.306	-74.597	1	7.8	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0026-A	13-SEP-2001	39.306	-74.597	2	7.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0028-A	17-JUL-2001	39.314	-74.629	1	3.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0030-C	29-AUG-2001	39.397	-74.39	1	2.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0032-A	17-JUL-2001	39.402	-74.718	1	2.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0034-A	29-AUG-2001	39.437	-74.381	1	0.5	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0036-A	08-AUG-2001	39.511	-74.297	1	4.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0036-A	07-SEP-2001	39.511	-74.297	1	6.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0038-A	19-JUL-2001	39.557	-74.48	1	7.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0040-A	20-JUL-2001	39.589	-74.24	1	2.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0042-A	25-JUL-2001	39.625	-74.236	1	0.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0042-A	27-JUL-2001	39.625	-74.236	2	1.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0042-A	31-OCT-2001	39.625	-74.236	3	1.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0044-A	10-AUG-2001	39.719	-74.173	1	0.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0046-A	24-JUL-2001	39.811	-74.168	1	1.5	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0046-A	31-OCT-2001	39.811	-74.168	2	2.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0048-A	24-JUL-2001	39.853	-74.102	1	1.4	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0050-A	23-JUL-2001	39.939	-74.091	1	1.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0050-A	31-OCT-2001	39.939	-74.091	2	1.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0052-A	23-JUL-2001	40.065	-74.133	1	1.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0054-A	12-JUL-2001	40.18	-74.044	1	2.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0056-A	12-JUL-2001	40.197	-74.037	1	1.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0058-C	27-AUG-2001	40.328	-74.01	1	1.8	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0060-A	19-SEP-2001	40.383	-73.98	1	2.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0060-A	30-OCT-2001	40.383	-73.98	2	2.1	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0062-A	15-OCT-2001	38.935	-74.98	1	11.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0064-A	13-SEP-2001	39.001	-74.957	1	1.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0066-B	13-SEP-2001	39.138	-74.968	1	3.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0068-A	23-AUG-2001	39.202	-75.041	1	2.5	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0070-B	06-OCT-2001	39.307	-75.329	1	5.8	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0072-A	23-AUG-2001	39.21	-75.099	1	2.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0074-A	09-OCT-2001	40.139	-74.732	1	5.4	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0076-A	08-OCT-2001	40.038	-74.989	1	5.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0078-A	10-OCT-2001	39.846	-75.265	1	12.1	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0080-A	15-OCT-2001	38.978	-75.1	1	11.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0082-A	20-SEP-2001	39.283	-75.242	1	2.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0084-A	22-AUG-2001	39.187	-74.912	1	1.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0086-A	20-SEP-2001	39.298	-75.18	1	0.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0088-A	20-AUG-2001	39.446	-75.411	1	0.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0090-A	19-SEP-2001	39.392	-75.041	1	3.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0102-A	05-OCT-2001	39.997	-74.113	1	1.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0104-A	04-OCT-2001	39.941	-74.179	1	1.8	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0106-A	04-OCT-2001	39.888	-74.111	1	1.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0108-A	08-OCT-2001	39.802	-74.174	1	0.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0110-A	08-OCT-2001	39.702	-74.179	1	0.5	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0112-A	10-OCT-2001	39.605	-74.261	1	2.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0114-A	11-OCT-2001	39.542	-74.309	1	0.8	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0116-A	11-OCT-2001	39.535	-74.377	1	1.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0118-A	12-OCT-2001	39.553	-74.454	1	3.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0120-A	18-OCT-2001	39.62	-74.63	1	1.8	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	NJ01-0122-A	18-OCT-2001	39.585	-74.538	1	0.8	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0003-A	07-OCT-2002	40.435	-74.038	1	6.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0013-A	05-SEP-2002	40.805	-74.14	1	5.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0023-A	26-SEP-2002	39.204	-74.655	1	3.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0033-A	26-SEP-2002	39.444	-74.454	1	1.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0043-A	04-SEP-2002	39.64	-74.205	1	1.5	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0053-A	27-AUG-2002	40.092	-74.078	1	2.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0073-A	05-AUG-2002	40.079	-74.87	1	14.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0075-A	06-AUG-2002	39.983	-75.067	1	14.4	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0077-A	06-AUG-2002	39.88	-75.179	1	14.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0079-A	06-AUG-2002	39.845	-75.338	1	12.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0081-A	30-JUL-2002	39.083	-75.183	1	13.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0200-A	06-SEP-2002	40.464	-74.251	1	2.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0203-A	06-SEP-2002	40.488	-74.422	1	2.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0205-A	10-OCT-2002	40.482	-74.036	1	5.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0206-A	10-OCT-2002	40.688	-74.126	1	10.5	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0208-A	05-SEP-2002	40.766	-74.157	1	3.5	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0211-A	07-OCT-2002	40.959	-73.905	1	13.4	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0213-A	25-SEP-2002	38.995	-74.828	1	1.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0214-A	25-SEP-2002	39.043	-74.772	1	3.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0216-A	25-SEP-2002	39.119	-74.722	1	3.1	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0219-A	24-SEP-2002	39.29	-74.659	1	3.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0221-A	11-SEP-2002	39.347	-74.709	1	4.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0222-A	24-SEP-2002	39.342	-74.478	1	5.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0224-A	11-SEP-2002	39.448	-74.729	1	0.8	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0227-A	23-SEP-2002	39.498	-74.334	1	1.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0229-A	03-SEP-2002	39.582	-74.536	1	1.5	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0230-A	15-AUG-2002	39.537	-74.334	1	1.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0232-A	03-SEP-2002	39.629	-74.643	1	0.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0235-A	04-SEP-2002	39.764	-74.108	1	8.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0237-C	28-AUG-2002	39.805	-74.102	1	1.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0238-A	28-AUG-2002	39.938	-74.11	1	1.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0240-A	27-AUG-2002	40.018	-74.073	1	1.8	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0243-A	29-AUG-2002	40.194	-74.035	1	0.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0245-C	16-AUG-2002	40.356	-74.078	1	0.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0246-A	16-AUG-2002	40.388	-74.015	1	0.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0249-A	29-JUL-2002	38.973	-74.981	1	5.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0249-A	30-JUL-2002	38.973	-74.981	2	6.1	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0251-A	30-JUL-2002	39.029	-75.081	1	7.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0251-A	31-JUL-2002	39.029	-75.081	2	7.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0253-A	31-JUL-2002	39.201	-75.22	1	5.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0255-A	03-OCT-2002	39.129	-74.922	1	2.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0257-A	19-SEP-2002	39.248	-75.207	1	3.5	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0259-A	19-SEP-2002	39.32	-75.333	1	5.4	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0260-A	14-OCT-2002	38.968	-74.961	1	1.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0261-A	14-OCT-2002	38.962	-74.924	1	3.1	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0262-A	03-OCT-2002	39.179	-74.836	1	1.5	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0264-A	18-SEP-2002	39.213	-75.104	1	1.8	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0266-A	19-SEP-2002	39.315	-75.288	1	1.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0268-A	01-OCT-2002	39.369	-75.035	1	0.5	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0270-A	01-OCT-2002	39.405	-75.232	1	0.8	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	NJ02-0272-C	17-SEP-2002	39.583	-75.493	1	8.8	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0008-A	28-OCT-2003	40.522	-73.97	1	6.5	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0018-A	23-OCT-2003	39.01	-74.842	1	1.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0028-A	21-OCT-2003	39.314	-74.629	1	1.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0038-A	29-OCT-2003	39.557	-74.48	1	7.8	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0048-A	04-SEP-2003	39.853	-74.102	1	1.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0058-A	14-AUG-2003	40.328	-74.01	1	0.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0074-A	04-AUG-2003	40.139	-74.732	1	6.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0076-A	04-AUG-2003	40.038	-74.989	1	5.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0078-A	05-AUG-2003	39.846	-75.265	1	10.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0080-A	29-JUL-2003	38.978	-75.1	1	11.4	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0201-A	17-SEP-2003	40.468	-74.158	1	4.5	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0204-A	28-OCT-2003	40.476	-74.214	1	4.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0207-A	16-SEP-2003	40.682	-74.058	1	2.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0209-A	15-SEP-2003	40.719	-74.11	1	1.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0210-A	15-SEP-2003	40.836	-74.029	1	0.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0212-A	23-OCT-2003	38.972	-74.846	1	5.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0217-A	30-OCT-2003	39.199	-74.688	1	2.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0218-A	24-OCT-2003	39.301	-74.773	1	0.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0220-A	30-OCT-2003	39.284	-74.582	1	1.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0225-A	21-OCT-2003	39.425	-74.714	1	1.8	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0234-A	05-SEP-2003	39.749	-74.187	1	1.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0236-B	05-SEP-2003	39.825	-74.16	1	1.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0239-A	04-SEP-2003	39.948	-74.102	1	2.1	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0241-A	31-OCT-2003	40.065	-74.133	1	1.1	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0242-A	19-AUG-2003	40.183	-74.052	1	0.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0244-A	19-AUG-2003	40.199	-74.043	1	1.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0247-A	20-AUG-2003	40.385	-73.981	1	1.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0248-A	28-JUL-2003	38.935	-74.979	1	11.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0252-A	09-OCT-2003	39.138	-74.967	1	3.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0254-A	17-OCT-2003	39.156	-75.034	1	3.1	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0256-A	08-OCT-2003	39.295	-75.316	1	2.5	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0258-A	17-OCT-2003	39.21	-75.098	1	2.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0263-A	08-OCT-2003	39.289	-75.207	1	3.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0269-B	08-OCT-2003	39.395	-75.412	1	7.4	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0271-A	20-OCT-2003	39.393	-75.04	1	3.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	NJ03-0273-A	07-OCT-2003	39.625	-75.487	1	1.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0003-A	30-JUN-2004	40.434	-74.038	1	5.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0013-A	17-AUG-2004	40.805	-74.14	1	6.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0023-A	27-SEP-2004	39.204	-74.655	1	1.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0033-A	15-SEP-2004	39.444	-74.454	1	1.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0043-A	28-JUL-2004	39.64	-74.205	1	1.8	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0053-A	20-JUL-2004	40.092	-74.078	1	1.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0073-A	09-AUG-2004	40.079	-74.87	1	14.1	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0077-A	11-AUG-2004	39.88	-75.179	1	8.5	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0215-A	23-SEP-2004	39.092	-74.796	1	0.4	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0223-B	17-SEP-2004	39.375	-74.409	1	7.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0226-B	15-SEP-2004	39.442	-74.348	1	1.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0228-A	18-AUG-2004	39.535	-74.268	1	1.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0231-A	27-JUL-2004	39.61	-74.218	1	2.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0233-A	27-JUL-2004	39.658	-74.219	1	0.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0250-A	22-SEP-2004	39.009	-74.959	1	4.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0252-A	21-SEP-2004	39.138	-74.967	1	4.4	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0265-A	21-SEP-2004	39.206	-74.922	1			
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0272-A	31-AUG-2004	39.583	-75.493	1	10.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0400-A	23-AUG-2004	40.485	-74.274	1	1.1	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0403-A	25-AUG-2004	40.487	-74.389	1	4.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0405-A	23-JUL-2004	40.478	-74.074	1	7.5	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0406-A	20-AUG-2004	40.656	-74.161	1	1.4	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0408-A	17-AUG-2004	40.735	-74.162	1	3.4	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0411-A	16-SEP-2004	40.954	-73.911	1	7.5	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0413-A	24-SEP-2004	39.009	-74.815	1	0.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0414-A	23-SEP-2004	39.06	-74.762	1	4.8	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0416-A	23-SEP-2004	39.115	-74.721	1	6.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0419-A	27-SEP-2004	39.307	-74.677	1	4.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0421-A	28-SEP-2004	39.366	-74.716	1	4.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0422-A	17-SEP-2004	39.363	-74.512	1	0.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0424-A	28-SEP-2004	39.444	-74.724	1	1.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0427-A	27-AUG-2004	39.521	-74.379	1	2.4	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0429-A	09-JUL-2004	39.568	-74.502	1	2.1	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0430-A	19-AUG-2004	39.575	-74.278	1	1.8	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0432-A	09-JUL-2004	39.62	-74.631	1	0.4	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0435-B	27-JUL-2004	39.721	-74.142	1	3.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0437-A	21-JUL-2004	39.818	-74.099	1	1.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0438-A	26-JUL-2004	39.944	-74.12	1	1.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0440-A	26-JUL-2004	40.04	-74.056	1	1.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0443-B	29-JUL-2004	40.194	-74.035	1	0.4	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0445-A	22-JUL-2004	40.339	-74.087	1	0.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0446-A	16-AUG-2004	40.38	-74.016	1	1.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0448-A	03-AUG-2004	38.975	-74.987	1	6.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0450-A	03-AUG-2004	39.112	-75.064	1	5.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0451-A	03-AUG-2004	39.197	-75.219	1	6.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0453-A	03-SEP-2004	39.134	-74.912	1	2.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0456-A	04-AUG-2004	39.313	-75.328	1	4.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0457-A	22-SEP-2004	38.966	-74.959	1	0.5	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0458-B	22-SEP-2004	38.966	-74.946	1	1.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0459-A	01-SEP-2004	39.282	-75.243	1	3.1	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0461-B	21-SEP-2004	39.176	-74.9	1	1.4	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0462-B	01-SEP-2004	39.299	-75.197	1	0.4	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0465-A	02-SEP-2004	39.429	-75.451	1	0.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0467-A	02-SEP-2004	39.387	-75.039	1	4.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0470-A	02-AUG-2004	38.96	-75.023	1	8.4	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0472-A	04-AUG-2004	39.261	-75.331	1	15.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	NJ04-0475-A	26-AUG-2004	40.133	-74.749	1	7.4	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2005	NJ05-0008-B	29-SEP-2005	40.652	-74.148	1		m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2005	NJ05-0011-A	05-OCT-2005	40.424	-74.053	1		m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2005	NJ05-0017-A	28-SEP-2005	40.498	-74.079	1		m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2005	NJ05-0020-A	28-SEP-2005	40.503	-73.989	1		m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2005	NJ05-0021-A	05-OCT-2005	40.464	-74.212	1		m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2005	NJ05-0025-B	05-OCT-2005	40.464	-74.122	1		m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2005	NJ05-0052-A	14-SEP-2005	39.885	-74.125	1		m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2005	NJ05-0054-B	16-SEP-2005	39.445	-74.383	1		m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2005	NJ05-0055-A	22-SEP-2005	40.461	-74.196	1		m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2005	NJ05-0056-A	20-SEP-2005	39.346	-74.53	1		m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2005	NJ05-0057-A	19-SEP-2005	39.584	-74.265	1		m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2005	NJ05-0058-A	19-SEP-2005	39.777	-74.154	1		m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2005	NJ05-0059-A	13-SEP-2005	39.505	-74.354	1		m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2005	NJ05-0060-A	22-SEP-2005	40.447	-74.074	1		m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2005	NJ05-021N-A	21-SEP-2005	40.358	-74.069	1		m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2005	NJ05-021T-A	21-SEP-2005	40.317	-73.995	1		m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0001-A	17-AUG-2006	39.942	-74.102	1	0.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0004-A	26-JUL-2006	39.626	-74.199	1	1.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0006-A	26-JUL-2006	39.565	-74.312	1	1.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0009-A	26-JUL-2006	39.568	-74.279	1	1.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0012-A	19-JUL-2006	39.847	-74.11	1	1.8	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0013-A	23-AUG-2006	39.365	-74.464	1	1.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0014-A	13-SEP-2006	40.939	-73.916	1	6.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0015-A	08-AUG-2006	39.536	-74.388	1	1.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0016-C	03-OCT-2006	40.494	-74.288	1	1.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0018-A	27-JUL-2006	39.523	-74.298	1	1.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0019-A	07-AUG-2006	39.277	-74.62	1	1.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0023-A	09-AUG-2006	39.043	-74.784	1	1.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0024-A	17-AUG-2006	40.003	-74.135	1	1.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0026-A	14-SEP-2006	40.476	-74.05	1	7.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0027-A	14-JUL-2006	39.5	-74.401	1	1.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0028-A	25-JUL-2006	39.438	-74.42	1	1.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0029-B	13-SEP-2006	40.695	-74.034	1	13.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0030-A	03-OCT-2006	40.473	-74.13	1	2.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0031-A	12-JUL-2006	39.787	-74.125	1	1.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0032-A	25-SEP-2006	40.43	-74.027	1	6.5	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0033-A	17-AUG-2006	40.063	-74.076	1	1.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0034-A	14-SEP-2006	40.486	-74.177	1	6.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0035-A	14-JUL-2006	39.496	-74.36	1	1.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0036-C	23-AUG-2006	39.29	-74.579	1	1.5	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0037-A	13-SEP-2006	40.679	-74.064	1	3.8	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0039-A	12-JUL-2006	39.73	-74.15	1	1.8	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0040-C	09-AUG-2006	38.966	-74.873	1	1.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0041-A	19-JUL-2006	39.867	-74.091	1	1.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0042-A	17-AUG-2006	39.947	-74.181	1	0.8	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0043-A	07-AUG-2006	39.294	-74.704	1	1.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0044-A	25-SEP-2006	40.415	-73.986	1	1.8	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0045-A	12-JUL-2006	39.666	-74.193	1	1.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0046-A	08-AUG-2006	39.612	-74.589	1	1.1	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0047-A	13-SEP-2006	40.787	-73.997	1	10.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0048-A	25-JUL-2006	39.45	-74.392	1	1.4	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0049-A	03-OCT-2006	40.503	-74.292	1	1.8	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0050-A	26-JUL-2006	39.595	-74.251	1	1.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0061-A	07-AUG-2006	39.366	-74.715	1	1.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0062-A	19-JUL-2006	39.852	-74.136	1	1.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0063-A	19-JUL-2006	39.904	-74.116	1	1.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0064-B	09-AUG-2006	39.037	-74.813	1	1.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0065-A	25-JUL-2006	39.473	-74.387	1	1.3	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0066-A	25-JUL-2006	39.396	-74.43	1	0.9	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0068-A	04-OCT-2006	40.381	-74.011	1	1.4	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0069-A	12-JUL-2006	39.616	-74.245	1	1.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2006	NJ06-0070-A	04-OCT-2006	40.357	-73.984	1	1.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0001-A	03-AUG-2000	40.776	-73.765	1	1.2	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0003-A	03-AUG-2000	40.785	-73.769	1	1.2	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0005-A	03-AUG-2000	40.835	-73.746	1	2.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0007-A	07-OCT-2000	40.856	-73.647	1	4.3	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0009-A	07-OCT-2000	40.871	-73.467	1	6.1	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0011-A	07-OCT-2000	40.882	-73.542	1	4.6	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0013-A	19-SEP-2000	40.922	-73.38	1	1.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0017-B	19-SEP-2000	40.927	-73.382	1	3.6	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0019-B	20-SEP-2000	40.955	-73.086	1	1.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0021-A	06-OCT-2000	41.126	-73.907	1	4.6	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0022-B	06-OCT-2000	41.279	-73.944	1	2.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0027-A	01-AUG-2000	40.506	-74.259	1	11.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0027-A	05-OCT-2000	40.506	-74.259	2	13.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0029-A	01-AUG-2000	40.573	-73.884	1	11.3	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0029-A	05-OCT-2000	40.573	-73.884	2	9.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0031-A	02-AUG-2000	40.644	-74.054	1	14.2	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0031-A	05-OCT-2000	40.644	-74.054	2	15.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0033-A	02-AUG-2000	40.765	-74.006	1	15.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0035-B	14-AUG-2000	40.802	-73.788	1	26.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0037-A	14-AUG-2000	40.806	-73.841	1	3.1	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0039-A	16-AUG-2000	40.594	-73.674	1	4.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0039-A	04-OCT-2000	40.594	-73.674	2	8.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0041-B	12-SEP-2000	40.618	-73.421	1	1.7	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0043-A	16-AUG-2000	40.621	-73.604	1	5.2	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0045-A	12-SEP-2000	40.68	-73.261	1	1.7	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0045-A	04-OCT-2000	40.68	-73.261	2	2.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0047-A	12-SEP-2000	40.689	-73.102	1	1.7	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0047-A	03-OCT-2000	40.689	-73.102	2	2.1	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0049-A	12-SEP-2000	40.708	-73.118	1	2.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0049-A	03-OCT-2000	40.708	-73.118	4	3.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0049-A	04-OCT-2000	40.708	-73.118	2	3.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0055-A	03-OCT-2000	40.86	-72.481	1	2.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0057-A	14-JUL-2000	40.931	-72.518	1	6.1	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0057-A	02-OCT-2000	40.931	-72.518	2	6.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0059-A	14-JUL-2000	41.0	-72.412	1	9.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0059-A	02-OCT-2000	41.0	-72.412	2	9.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0061-A	13-JUL-2000	41.059	-72.148	1	7.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0063-A	12-JUL-2000	41.05	-71.916	1	2.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0065-A	13-JUL-2000	41.108	-72.193	1	9.6	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2000	NY00-0067-A	12-JUL-2000	41.066	-71.921	1	2.6	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	NY00-0069-A	07-AUG-2000	40.935	-73.6	1	15.2	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	NY00-0071-A	08-AUG-2000	40.961	-73.476	1	17.3	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	NY00-0073-A	21-JUL-2000	40.952	-73.332	1	16.1	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	NY00-0075-A	17-AUG-2000	41.055	-73.08	1	24.2	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	NY00-0079-A	30-AUG-2000	41.004	-72.768	1	25.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	NY00-0081-A	15-AUG-2000	41.098	-72.45	1	18.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	NY00-0083-A	07-AUG-2000	40.873	-73.734	1	33.3	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	NY00-0085-A	10-JUL-2000	40.956	-73.58	1	18.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	NY00-0087-A	02-AUG-2000	41.026	-72.913	1	40.0	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	NY00-0091-A	04-AUG-2000	41.262	-72.009	1	3.5	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	NY00-0093-B	14-SEP-2000	40.996	-73.032	1	22.9	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	NY00-0095-A	12-SEP-2000	41.044	-72.601	1	21.6	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	NY00-0097-A	14-SEP-2000	41.057	-72.927	1	32.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	NY00-0099-A	11-SEP-2000	41.084	-72.538	1	24.2	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	NY00-0101-A	13-SEP-2000	41.09	-72.794	1	31.6	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	NY00-0103-A	11-SEP-2000	41.109	-72.617	1	25.8	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	NY00-0105-A	13-SEP-2000	41.129	-72.697	1	30.4	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	NY00-0107-A	11-SEP-2000	41.143	-72.626	1	28.2	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	NY00-0109-A	21-SEP-2000	40.93	-73.204	1	15.4	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	NY00-0111-A	21-SEP-2000	40.968	-73.396	1	14.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2000	NY00-0113-A	14-SEP-2000	41.001	-72.973	1	18.3	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0002-A	06-AUG-2001	40.797	-73.772	1	3.7	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0002-A	23-AUG-2001	40.797	-73.772	2	2.7	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0004-B	06-AUG-2001	40.833	-73.655	1	6.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0006-A	06-AUG-2001	40.833	-73.717	1	2.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0006-A	23-AUG-2001	40.833	-73.717	2	2.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0008-A	08-AUG-2001	40.877	-73.54	1	3.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0012-B	07-AUG-2001	40.896	-73.498	1	4.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0012-B	08-AUG-2001	40.896	-73.498	2	5.2	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0014-A	07-AUG-2001	40.918	-73.364	1	3.7	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0014-A	09-AUG-2001	40.918	-73.364	2	4.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0016-A	08-AUG-2001	40.919	-73.161	1	1.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0016-A	09-AUG-2001	40.919	-73.161	2	3.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0018-A	09-AUG-2001	40.968	-73.087	1	5.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0018-A	10-AUG-2001	40.968	-73.087	2	5.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0020-B	10-AUG-2001	40.97	-73.084	1	5.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0023-A	31-JUL-2001	41.931	-73.955	1	8.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0024-A	01-AUG-2001	42.656	-73.74	1	7.6	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0025-A	01-AUG-2001	42.745	-73.687	1	6.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0026-A	16-AUG-2001	40.501	-74.149	1	7.3	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0026-A	24-AUG-2001	40.501	-74.149	2	7.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0028-A	26-JUL-2001	40.568	-73.983	1	5.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0028-A	21-AUG-2001	40.568	-73.983	2	4.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0030-A	24-AUG-2001	40.638	-74.195	1	12.2	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0032-A	26-JUL-2001	40.627	-73.882	1	9.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0032-A	21-AUG-2001	40.627	-73.882	2	11.3	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0034-A	22-AUG-2001	40.788	-73.935	1	5.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0036-B	22-AUG-2001	40.878	-73.924	1	6.7	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0038-A	30-JUL-2001	40.915	-73.916	1	14.3	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0040-A	25-JUL-2001	40.621	-73.508	1	3.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0042-A	24-JUL-2001	40.634	-73.254	1	7.3	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0042-A	30-JUL-2001	40.634	-73.254	2	2.1	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0044-A	25-JUL-2001	40.649	-73.476	1	3.7	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0046-A	23-JUL-2001	40.682	-73.205	1	1.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0046-A	30-JUL-2001	40.682	-73.205	2	1.1	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0048-A	23-JUL-2001	40.708	-73.236	1	2.1	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0048-A	30-JUL-2001	40.708	-73.236	2	1.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0050-A	23-JUL-2001	40.741	-72.998	1	2.3	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0050-A	31-JUL-2001	40.741	-72.998	1	2.1	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0052-A	23-JUL-2001	40.792	-72.718	1	1.7	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0052-A	31-JUL-2001	40.792	-72.718	2	1.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0054-B	20-JUL-2001	40.848	-72.543	1	1.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0054-B	01-AUG-2001	40.848	-72.543	1	1.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0056-A	20-JUL-2001	40.929	-72.607	1	2.1	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0056-A	24-JUL-2001	40.929	-72.607	2	2.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0058-A	16-JUL-2001	40.96	-72.424	1	8.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0058-A	17-JUL-2001	40.96	-72.424	2	6.7	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0060-A	18-JUL-2001	41.039	-72.33	1	8.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0060-A	23-JUL-2001	41.039	-72.33	2	8.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0060-B	18-JUL-2001	41.036	-72.245	2	3.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0060-B	23-JUL-2001	41.036	-72.245	1	3.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0062-B	19-JUL-2001	41.07	-72.035	1	12.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0062-B	25-JUL-2001	41.07	-72.035	2	14.6	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0064-C	24-JUL-2001	41.091	-72.353	1	5.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0066-A	19-JUL-2001	41.077	-72.076	1	7.3	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0066-A	25-JUL-2001	41.077	-72.076	2	7.3	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0066-C	19-JUL-2001	41.08	-72.103	2	5.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0066-C	25-JUL-2001	41.08	-72.103	1	5.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0068-A	19-JUL-2001	41.173	-72.163	1	10.3	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2001	NY01-0068-A	26-JUL-2001	41.173	-72.163	2	11.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	NY01-0070-A	25-JUL-2001	40.938	-73.519	1	10.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	NY01-0072-A	21-AUG-2001	40.95	-73.425	1	11.2	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	NY01-0074-A	01-AUG-2001	40.992	-73.218	1	25.6	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	NY01-0076-A	01-AUG-2001	40.994	-73.042	1	22.1	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	NY01-0077-A	22-AUG-2001	40.981	-72.918	1	10.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	NY01-0078-A	29-AUG-2001	41.078	-72.833	1	29.1	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	NY01-0079-A	29-AUG-2001	41.004	-72.768	1	25.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	NY01-0080-A	08-AUG-2001	41.004	-72.651	1	19.8	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	NY01-0082-A	11-JUL-2001	40.931	-73.221	1	14.2	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	NY01-0084-A	10-JUL-2001	40.918	-73.642	1	17.8	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	NY01-0086-A	01-AUG-2001	41.018	-73.144	1	39.8	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	NY01-0088-A	09-JUL-2001	41.138	-72.655	1	26.1	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	NY01-0089-A	29-AUG-2001	41.182	-72.457	1	21.8	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2001	NY01-0090-A	09-AUG-2001	41.237	-72.053	1	73.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0001-A	03-MAY-2002	40.776	-73.765	1	2.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0001-A	10-SEP-2002	40.776	-73.765	2	2.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0003-A	03-MAY-2002	40.785	-73.769	1	3.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0005-A	02-MAY-2002	40.835	-73.746	1	4.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0006-A	12-AUG-2002	40.833	-73.717	1	2.7	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0006-A	09-SEP-2002	40.833	-73.717	2	2.1	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0007-A	06-MAY-2002	40.856	-73.647	1	7.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0007-A	10-SEP-2002	40.856	-73.647	2	7.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0009-A	07-MAY-2002	40.871	-73.467	1	6.1	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0011-A	07-MAY-2002	40.882	-73.542	1	5.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0011-A	13-SEP-2002	40.882	-73.542	2	5.6	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0013-B	08-MAY-2002	40.923	-73.422	1	7.3	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0013-B	13-SEP-2002	40.923	-73.422	2	8.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0016-A	20-AUG-2002	40.919	-73.161	1	4.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0016-A	21-AUG-2002	40.919	-73.161	2	3.7	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0017-A	08-MAY-2002	40.927	-73.381	1	5.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0017-A	12-SEP-2002	40.927	-73.381	2	6.3	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0019-B	09-MAY-2002	40.955	-73.086	1	9.1	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0019-B	11-SEP-2002	40.955	-73.086	2	8.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0029-A	14-AUG-2002	40.573	-73.884	1	10.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0029-A	03-SEP-2002	40.573	-73.884	2	10.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0044-A	30-AUG-2002	40.649	-73.476	1	3.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0052-A	17-JUL-2002	40.792	-72.718	1	1.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0052-A	05-AUG-2002	40.792	-72.718	2	2.1	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0057-A	10-JUL-2002	40.931	-72.518	1	6.3	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0057-A	31-JUL-2002	40.931	-72.518	2	6.7	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0201-A	12-AUG-2002	40.799	-73.777	1	7.6	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0201-A	10-SEP-2002	40.799	-73.777	2	3.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0204-A	12-AUG-2002	40.843	-73.734	1	4.6	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0204-A	09-SEP-2002	40.843	-73.734	2	5.1	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0207-B	16-AUG-2002	40.869	-73.472	1	1.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0207-B	13-SEP-2002	40.869	-73.472	2	4.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0210-A	16-AUG-2002	40.882	-73.474	1	6.3	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0210-A	13-SEP-2002	40.882	-73.474	2	4.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0216-A	19-AUG-2002	40.965	-73.082	1	10.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0216-A	11-SEP-2002	40.965	-73.082	2	7.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0223-A	15-AUG-2002	40.492	-74.253	1	13.7	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0223-A	04-SEP-2002	40.492	-74.253	2	12.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0226-A	13-AUG-2002	40.521	-74.01	1	11.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0226-A	04-SEP-2002	40.521	-74.01	2	10.1	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0229-A	13-AUG-2002	40.544	-74.047	1	10.1	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0229-A	04-SEP-2002	40.544	-74.047	2	10.1	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0232-A	13-AUG-2002	40.644	-74.053	1	15.2	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0232-A	05-SEP-2002	40.644	-74.053	2	15.1	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0235-A	14-AUG-2002	40.646	-73.82	1	8.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0235-A	03-SEP-2002	40.646	-73.82	2	7.7	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0237-A	14-AUG-2002	40.664	-74.031	1	4.6	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0237-A	05-SEP-2002	40.664	-74.031	2	4.6	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0239-A	14-AUG-2002	40.659	-73.839	1	11.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0242-A	15-AUG-2002	40.796	-73.794	1	10.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0242-A	09-SEP-2002	40.796	-73.794	2	10.6	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0243-A	15-AUG-2002	40.836	-73.959	1	11.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0243-A	06-SEP-2002	40.836	-73.959	2	10.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0248-A	28-AUG-2002	40.614	-73.449	1	4.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0250-B	29-AUG-2002	40.623	-73.611	1	3.6	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0251-B	18-JUL-2002	40.673	-73.329	1	3.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0251-B	06-AUG-2002	40.673	-73.329	2	2.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0253-B	18-JUL-2002	40.689	-73.074	1	2.2	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0253-B	05-AUG-2002	40.689	-73.074	2	3.7	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0258-A	17-JUL-2002	40.809	-72.725	1	0.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0258-A	05-AUG-2002	40.809	-72.725	2	2.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0260-A	17-JUL-2002	40.878	-72.474	1	2.3	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-0260-A	01-AUG-2002	40.878	-72.474	2	2.8	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	NY02-0275-A	18-SEP-2002	41.04	-72.649	1	22.6	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	NY02-0276-A	30-SEP-2002	41.056	-72.928	1	31.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	NY02-0277-A	23-SEP-2002	41.063	-72.834	1	30.5	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	NY02-0278-A	19-SEP-2002	41.077	-72.76	1	29.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	NY02-0279-A	18-SEP-2002	41.089	-72.755	1	28.4	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	NY02-0280-A	18-SEP-2002	41.115	-72.568	1	25.3	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	NY02-0281-A	20-SEP-2002	41.136	-72.675	1	27.4	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	NY02-0282-A	17-SEP-2002	41.132	-72.495	1	28.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	NY02-0283-A	17-SEP-2002	41.15	-72.495	1	41.2	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	NY02-0284-A	01-OCT-2002	40.924	-73.591	1	12.5	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	NY02-0285-A	02-OCT-2002	40.935	-73.68	1	12.5	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	NY02-0286-A	19-SEP-2002	40.978	-72.745	1	10.4	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2002	NY02-0287-A	30-SEP-2002	40.993	-72.999	1	18.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-1001-A	12-JUL-2002	41.152	-72.243	1	3.7	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-1001-A	25-JUL-2002	41.152	-72.243	2	4.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-1002-B	16-JUL-2002	41.105	-72.145	1	8.3	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-1002-B	25-JUL-2002	41.105	-72.145	2	9.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-1003-A	22-JUL-2002	41.089	-72.019	1	15.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-1003-A	29-JUL-2002	41.089	-72.019	2	17.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-1004-B	22-JUL-2002	41.051	-72.032	1	0.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-1004-B	29-JUL-2002	41.051	-72.032	2	8.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-1006-A	08-JUL-2002	41.126	-72.27	1	3.3	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-1006-A	25-JUL-2002	41.126	-72.27	2	6.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-1007-A	08-JUL-2002	41.133	-72.318	1	5.3	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-1007-A	30-JUL-2002	41.133	-72.318	2	5.6	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-1011-A	12-JUL-2002	41.085	-72.211	1	11.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-1011-A	23-JUL-2002	41.085	-72.211	2	11.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-1015-A	09-JUL-2002	41.076	-72.389	1	10.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-1015-A	30-JUL-2002	41.076	-72.389	2	14.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-1016-A	09-JUL-2002	41.052	-72.309	1	3.3	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-1016-A	26-JUL-2002	41.052	-72.309	2	6.6	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-1017-A	15-JUL-2002	40.998	-72.1	1	3.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-1017-A	23-JUL-2002	40.998	-72.1	2	4.2	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-1019-B	15-JUL-2002	41.041	-72.199	1	7.7	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-1019-B	23-JUL-2002	41.041	-72.199	2	8.2	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-1020-A	16-JUL-2002	41.002	-72.183	1	2.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-1021-A	09-JUL-2002	41.021	-72.333	1	4.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-1021-A	26-JUL-2002	41.021	-72.333	2	9.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-1022-A	10-JUL-2002	41.027	-72.406	1	2.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-1022-A	24-JUL-2002	41.027	-72.406	2	3.6	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-1025-A	10-JUL-2002	40.976	-72.528	1	1.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-1025-A	24-JUL-2002	40.976	-72.528	2	4.1	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-1026-A	11-JUL-2002	40.951	-72.417	1	1.7	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-1026-A	31-JUL-2002	40.951	-72.417	2	5.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-1027-A	11-JUL-2002	40.927	-72.471	1	7.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-1027-A	31-JUL-2002	40.927	-72.471	2	7.7	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-1030-A	11-JUL-2002	40.913	-72.59	1	1.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2002	NY02-1030-A	01-AUG-2002	40.913	-72.59	2	5.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2003	NY03-0072-A	20-AUG-2003	40.95	-73.425	1	11.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2003	NY03-0074-A	21-AUG-2003	40.992	-73.218	1	24.3	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2003	NY03-0075-A	25-JUL-2003	41.055	-73.08	1	25.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0084-A	02-MAY-2003	40.918	-73.642	1	17.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0084-A	11-AUG-2003	40.918	-73.642	3	18.2	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0084-A	12-AUG-2003	40.918	-73.642	4	17.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0084-A	14-AUG-2003	40.918	-73.642	5	16.9	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2003	NY03-0084-X	28-JUL-2003	40.918	-73.642	2	17.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2003	NY03-0088-A	24-JUL-2003	41.138	-72.655	1	27.2	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2003	NY03-0088-A	19-AUG-2003	41.138	-72.655	2	26.2	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2003	NY03-0089-A	27-AUG-2003	41.182	-72.457	1	29.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0202-A	02-MAY-2003	40.826	-73.731	1	5.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0202-B	04-AUG-2003	40.83	-73.725	2	4.3	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0202-B	15-AUG-2003	40.83	-73.725	3	4.7	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0205-A	01-MAY-2003	40.855	-73.647	1	8.6	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0205-C	11-AUG-2003	40.856	-73.646	2	4.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0205-C	14-AUG-2003	40.856	-73.646	3	8.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0211-A	05-MAY-2003	40.908	-73.406	1	6.7	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0211-A	12-AUG-2003	40.908	-73.406	2	7.2	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0211-A	19-AUG-2003	40.908	-73.406	3	8.6	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0214-A	05-MAY-2003	40.924	-73.372	1	4.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0214-A	12-AUG-2003	40.924	-73.372	2	5.3	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0214-A	19-AUG-2003	40.924	-73.372	3	4.3	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0217-A	07-MAY-2003	40.97	-73.084	1	9.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0217-A	13-AUG-2003	40.97	-73.084	2	7.2	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0217-A	19-AUG-2003	40.97	-73.084	3	8.6	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0224-A	06-AUG-2003	40.517	-74.169	1	4.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0224-A	07-AUG-2003	40.517	-74.169	2	4.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0227-A	06-AUG-2003	40.58	-74.21	1	13.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0227-A	07-AUG-2003	40.58	-74.21	2	11.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0230-A	05-AUG-2003	40.561	-73.958	1	7.6	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0230-A	06-AUG-2003	40.561	-73.958	2	5.6	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0233-A	05-AUG-2003	40.6	-74.031	1	15.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0233-A	06-AUG-2003	40.6	-74.031	2	9.3	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0236-A	05-AUG-2003	40.631	-73.742	1	3.3	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0240-A	06-AUG-2003	40.747	-73.96	1	12.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0240-A	08-AUG-2003	40.747	-73.96	2	11.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0244-C	04-AUG-2003	40.801	-73.818	1	12.2	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0244-C	08-AUG-2003	40.801	-73.818	2	12.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0249-A	16-JUL-2003	40.631	-73.248	1	8.3	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0249-A	05-AUG-2003	40.631	-73.248	2	8.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0252-B	14-JUL-2003	40.692	-73.168	1	3.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0252-B	05-AUG-2003	40.692	-73.168	2	2.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0255-A	14-JUL-2003	40.704	-73.123	1	3.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0255-A	05-AUG-2003	40.704	-73.123	2	2.7	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0259-A	10-JUL-2003	40.847	-72.543	1	1.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0259-A	04-AUG-2003	40.847	-72.543	2	1.7	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0261-B	10-JUL-2003	40.933	-72.601	1	3.3	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0263-A	09-JUL-2003	41.009	-72.409	1	4.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0263-A	30-JUL-2003	41.009	-72.409	2	11.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0265-A	09-JUL-2003	41.043	-72.08	1	5.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0265-A	01-AUG-2003	41.043	-72.08	2	5.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0267-B	31-JUL-2003	41.052	-71.917	1	2.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0268-A	08-JUL-2003	41.105	-72.312	1	5.2	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0268-A	30-JUL-2003	41.105	-72.312	2	5.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0269-A	08-JUL-2003	41.12	-72.282	1	1.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0269-A	01-AUG-2003	41.12	-72.282	2	6.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2003	NY03-0271-C	31-JUL-2003	41.063	-71.923	1	2.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2003	NY03-0291-A	16-SEP-2003	41.036	-72.701	1	27.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2003	NY03-0292-A	11-SEP-2003	41.058	-72.709	1	26.5	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2003	NY03-0293-A	29-SEP-2003	40.931	-73.544	1	11.6	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2003	NY03-0294-A	16-SEP-2003	40.976	-72.746	1	9.1	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2003	NY03-0295-A	24-SEP-2003	40.983	-72.948	1	10.1	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2004	NY04-0070-A	03-SEP-2004	40.938	-73.519	1	11.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2004	NY04-0072-A	03-SEP-2004	40.95	-73.425	1	11.4	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2004	NY04-0075-A	07-SEP-2004	41.055	-73.08	1	24.8	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2004	NY04-0080-A	19-JUL-2004	41.004	-72.651	1	20.7	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2004	NY04-0082-A	21-JUL-2004	40.931	-73.221	1	15.2	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0083-A	02-AUG-2004	40.873	-73.734	1	35.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0083-A	08-SEP-2004	40.873	-73.734	2	12.8	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2004	NY04-0083-X	20-JUL-2004	40.873	-73.734	1	34.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2004	NY04-0087-A	19-AUG-2004	41.026	-72.913	1	40.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0200-A	14-JUL-2004	40.775	-73.76	1	3.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0200-A	09-SEP-2004	40.775	-73.76	2	4.1	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0206-A	15-JUL-2004	40.879	-73.516	2	5.3	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0206-A	13-SEP-2004	40.879	-73.516	3	3.2	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0209-B	15-JUL-2004	40.884	-73.541	1	6.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0209-B	13-SEP-2004	40.884	-73.541	2	8.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0212-B	15-JUL-2004	40.918	-73.358	1	4.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0212-B	10-SEP-2004	40.918	-73.358	2	5.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0218-A	19-JUL-2004	41.075	-73.892	1	5.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0219-A	19-JUL-2004	41.186	-73.919	1	4.2	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0220-A	20-JUL-2004	42.096	-73.927	1	8.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0221-A	21-JUL-2004	42.505	-73.777	1	12.3	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0222-A	21-JUL-2004	42.729	-73.696	1	6.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0225-A	12-JUL-2004	40.522	-74.107	1	5.1	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0225-A	03-AUG-2004	40.522	-74.107	2	6.7	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0228-C	12-JUL-2004	40.546	-74.103	1	2.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0228-C	03-AUG-2004	40.546	-74.103	2	3.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0231-A	09-JUL-2004	40.609	-74.2	1	3.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0231-B	04-AUG-2004	40.642	-74.155	2	4.3	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0234-A	12-JUL-2004	40.608	-73.882	1	14.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0234-A	03-AUG-2004	40.608	-73.882	2	12.2	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0238-B	04-AUG-2004	40.708	-73.987	1	16.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0241-B	13-JUL-2004	40.793	-73.876	1	14.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0241-C	02-AUG-2004	40.786	-73.921	2	8.2	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0245-A	13-JUL-2004	40.875	-73.916	1	8.7	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0245-A	04-AUG-2004	40.875	-73.916	2	12.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0246-B	08-JUL-2004	40.611	-73.631	1	6.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0254-A	07-JUL-2004	40.71	-73.232	1	1.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0254-A	15-SEP-2004	40.71	-73.232	2	2.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0256-A	07-JUL-2004	40.741	-73.015	1	1.7	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0256-A	14-SEP-2004	40.741	-73.015	2	2.7	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0262-A	27-JUL-2004	40.949	-72.437	2	2.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0262-B	27-JUL-2004	40.971	-72.393	1	8.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0264-A	26-JUL-2004	41.054	-72.239	1	6.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0264-A	27-JUL-2004	41.054	-72.239	2	4.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0266-A	26-JUL-2004	41.054	-71.999	1	16.2	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0266-A	28-JUL-2004	41.054	-71.999	2	15.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0270-B	26-JUL-2004	41.088	-72.06	1	8.2	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0270-B	28-JUL-2004	41.088	-72.06	2	7.6	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0272-A	23-JUL-2004	41.167	-72.156	1	13.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2004	NY04-0272-A	29-JUL-2004	41.167	-72.156	2	14.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2004	NY04-0284-A	30-SEP-2004	40.925	-73.593	1	14.9	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2004	NY04-0401-A	15-SEP-2004	41.019	-72.808	1	36.0	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2004	NY04-0405-A	13-SEP-2004	41.121	-72.518	1	30.8	m	
National Coastal Assessment-Northeast/Connecticut Dept. of Environmental Protection	2004	NY04-0409-A	16-SEP-2004	40.992	-72.818	1	5.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0001-A	19-JUL-2005	40.649	-73.177	1	3.3	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0001-A	02-AUG-2005	40.649	-73.177	2	7.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0002-B	14-JUL-2005	40.594	-73.873	1	4.1	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0002-B	09-AUG-2005	40.594	-73.873	2	10.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0003-A	12-JUL-2005	41.237	-73.969	1	4.3	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0004-B	11-JUL-2005	40.926	-73.383	1	3.2	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0005-A	27-JUL-2005	41.025	-72.358	1	12.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0005-A	14-SEP-2005	41.025	-72.358	2	7.2	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0006-A	26-JUL-2005	41.087	-72.044	1	12.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0006-A	13-SEP-2005	41.087	-72.044	2	10.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0007-B	25-JUL-2005	40.897	-72.491	1	1.1	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0007-B	14-SEP-2005	40.897	-72.491	2	8.1	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0008-A	26-JUL-2005	41.096	-72.17	1	9.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0008-A	12-SEP-2005	41.096	-72.17	2	10.1	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0009-B	19-JUL-2005	40.695	-73.156	1	3.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0009-B	02-AUG-2005	40.695	-73.156	2	2.6	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0010-B	09-AUG-2005	40.629	-73.749	2	2.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0010-C	14-JUL-2005	40.632	-73.807	1	10.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0011-A	18-JUL-2005	40.619	-73.498	1	2.2	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0012-A	20-JUL-2005	40.717	-72.993	1	3.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0012-A	01-AUG-2005	40.717	-72.993	2	2.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0013-C	03-AUG-2005	40.855	-72.478	1	1.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0013-C	15-SEP-2005	40.855	-72.478	2	2.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0014-A	26-JUL-2005	41.07	-72.176	1	12.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0014-A	13-SEP-2005	41.07	-72.176	2	11.1	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0015-A	14-JUL-2005	40.514	-74.163	1	6.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0015-A	09-AUG-2005	40.514	-74.163	2	5.3	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0016-A	26-JUL-2005	41.035	-72.021	1	12.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0016-A	13-SEP-2005	41.035	-72.021	2	10.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0017-A	13-JUL-2005	40.538	-73.958	1	9.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0017-A	09-AUG-2005	40.538	-73.958	2	8.6	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0018-A	26-JUL-2005	41.022	-72.07	1	7.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0019-A	25-JUL-2005	40.973	-72.52	1	1.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0019-A	15-SEP-2005	40.973	-72.52	2	6.6	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0020-A	27-JUL-2005	41.079	-72.311	1	2.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0020-C	13-SEP-2005	41.094	-72.287	2	5.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0021-A	08-AUG-2005	40.699	-74.02	2	9.2	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0021-B	13-JUL-2005	40.678	-74.036	1	10.1	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0022-A	25-JUL-2005	40.961	-72.4	1	1.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0022-A	14-SEP-2005	40.961	-72.4	2	8.6	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0023-A	12-JUL-2005	40.801	-73.828	1	7.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0024-A	19-JUL-2005	40.702	-73.047	1	3.6	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0024-A	01-AUG-2005	40.702	-73.047	2	3.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0025-A	13-JUL-2005	40.605	-74.033	1	10.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2005	NY05-0025-A	08-AUG-2005	40.605	-74.033	2	4.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0026-A	09-AUG-2006	41.543	-73.985	1	11.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0026-A	10-AUG-2006	41.543	-73.985	2	8.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0027-A	08-AUG-2006	40.533	-74.069	1	6.1	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0027-A	14-AUG-2006	40.533	-74.069	2	4.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0028-A	07-JUL-2006	40.932	-72.516	1	7.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0028-A	17-JUL-2006	40.932	-72.516	1	7.3	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0029-A	06-JUL-2006	41.068	-72.248	1	5.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0029-A	12-SEP-2006	41.068	-72.248	2	12.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0030-A	07-AUG-2006	40.574	-74.025	1	10.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0030-A	14-AUG-2006	40.574	-74.025	2	10.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0031-A	07-JUL-2006	41.022	-72.375	1	7.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0031-A	11-SEP-2006	41.022	-72.375	2	7.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0032-C	13-JUL-2006	40.673	-73.32	1	1.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0032-C	28-JUL-2006	40.673	-73.32	2	1.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0033-A	12-JUL-2006	40.786	-72.724	1	1.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0034-A	07-AUG-2006	40.564	-73.923	1	6.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0034-A	15-AUG-2006	40.564	-73.923	2	12.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0035-C	06-JUL-2006	41.007	-72.089	1	2.7	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0035-C	12-SEP-2006	41.007	-72.089	2	3.7	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0036-B	07-JUL-2006	40.925	-72.609	1	1.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0036-B	18-JUL-2006	40.925	-72.609	2	3.1	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0037-A	05-JUL-2006	41.127	-72.232	1	11.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0037-A	13-SEP-2006	41.127	-72.232	2	11.2	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0038-A	09-AUG-2006	41.087	-73.908	1	4.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0038-A	10-AUG-2006	41.087	-73.908	2	4.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0039-B	06-JUL-2006	41.081	-72.376	1	1.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0039-B	11-SEP-2006	41.081	-72.376	2	4.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0040-A	11-AUG-2006	40.798	-73.766	1	2.5	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0041-A	12-JUL-2006	40.717	-73.053	1	2.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0041-A	26-JUL-2006	40.717	-73.053	1	3.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0042-A	12-JUL-2006	40.676	-73.104	1	1.7	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0042-A	26-JUL-2006	40.676	-73.104	2	2.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0043-A	07-AUG-2006	40.633	-73.802	1	10.1	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0043-A	15-AUG-2006	40.633	-73.802	2	5.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0044-B	01-AUG-2006	40.628	-73.493	1	6.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0044-B	03-AUG-2006	40.628	-73.493	2	3.0	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0045-B	12-JUL-2006	40.755	-72.908	1		m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0045-B	27-JUL-2006	40.755	-72.908	2	2.2	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0046-A	06-JUL-2006	41.004	-72.277	1	3.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0046-A	11-SEP-2006	41.004	-72.277	2	4.3	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0047-A	06-JUL-2006	41.044	-72.133	1	4.7	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0047-A	12-SEP-2006	41.044	-72.133	2	8.9	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0048-A	08-AUG-2006	40.491	-74.241	1	5.8	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0048-A	14-AUG-2006	40.491	-74.241	2	3.4	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0049-A	05-JUL-2006	41.128	-72.267	1	3.6	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0049-A	13-SEP-2006	41.128	-72.267	2	8.1	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0050-A	12-JUL-2006	40.67	-73.215	1	3.7	m	
National Coastal Assessment-Northeast/MSRC/Stonybrook U./Suffolk Co. Dept. HS/NYC DEP/Hempstead	2006	NY06-0050-A	28-JUL-2006	40.67	-73.215	2	2.4	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2000	PA00-0003-C	27-SEP-2000	39.954	-75.181	1	4.7	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	PA01-0002-A	09-OCT-2001	39.951	-75.137	1	14.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2001	PA01-0004-A	26-SEP-2001	39.913	-75.205	1	12.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2002	PA02-0201-B	16-SEP-2002	39.962	-75.182	1	8.0	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	PA03-0002-A	05-AUG-2003	39.951	-75.137	1	15.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2003	PA03-0200-A	03-OCT-2003	39.928	-75.212	1	4.6	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	PA04-0400-C	10-AUG-2004	39.928	-75.211	1	5.1	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	PA04-0402-A	11-AUG-2004	39.812	-75.397	1	15.2	m	
National Coastal Assessment-Northeast/New Jersey Marine Sciences Consortium	2004	PA04-0404-C	10-AUG-2004	39.921	-75.133	1	17.2	m	
R-EMAP Region 2 1993-94	1993	RB001	12-AUG-1993	40.581	-74.035	1	20.7	m	
R-EMAP Region 2 1998	1998	RB001	01-JUL-1998	40.58	-74.034	1			
R-EMAP Region 2 1998	1998	RB001	04-JUL-1998	40.58	-74.034	2	21.0	m	
R-EMAP Region 2 1993-94	1993	RB002	12-AUG-1993	40.571	-74.08	1	4.0	m	
R-EMAP Region 2 1998	1998	RB002	01-JUL-1998	40.571	-74.081	1			
R-EMAP Region 2 1998	1998	RB002	06-JUL-1998	40.571	-74.081	2	3.5	m	
R-EMAP Region 2 1993-94	1993	RB007	12-AUG-1993	40.547	-74.085	1	6.4	m	
R-EMAP Region 2 1998	1998	RB007	01-JUL-1998	40.546	-74.085	1			
R-EMAP Region 2 1998	1998	RB007	06-JUL-1998	40.546	-74.085	2	5.2	m	
R-EMAP Region 2 1993-94	1993	RB010	15-AUG-1993	40.538	-74.064	1	5.8	m	
R-EMAP Region 2 1998	1998	RB010	01-JUL-1998	40.538	-74.064	1			
R-EMAP Region 2 1998	1998	RB010	04-JUL-1998	40.538	-74.064	2	5.8	m	
R-EMAP Region 2 1993-94	1993	RB011	15-AUG-1993	40.535	-74.081	1	4.9	m	
R-EMAP Region 2 1998	1998	RB011	01-JUL-1998	40.535	-74.082	1			
R-EMAP Region 2 1998	1998	RB011	04-JUL-1998	40.535	-74.082	2	5.8	m	
R-EMAP Region 2 1993-94	1993	RB012	15-AUG-1993	40.533	-74.118	1	2.7	m	
R-EMAP Region 2 1998	1998	RB012	01-JUL-1998	40.534	-74.118	1			
R-EMAP Region 2 1998	1998	RB012	25-JUL-1998	40.534	-74.118	2	3.0	m	
R-EMAP Region 2 1993-94	1993	RB016	15-AUG-1993	40.507	-74.151	1	6.4	m	
R-EMAP Region 2 1998	1998	RB016	01-JUL-1998	40.507	-74.151	1			
R-EMAP Region 2 1998	1998	RB016	23-JUL-1998	40.507	-74.151	2	6.7	m	
R-EMAP Region 2 1993-94	1993	RB019	02-SEP-1993	40.495	-74.212	1	5.5	m	
R-EMAP Region 2 1998	1998	RB019	01-JUL-1998	40.496	-74.212	1			
R-EMAP Region 2 1998	1998	RB019	24-JUL-1998	40.496	-74.212	2	4.9	m	
R-EMAP Region 2 1993-94	1993	RB024	17-AUG-1993	40.474	-74.048	1	7.6	m	
R-EMAP Region 2 1998	1998	RB024	01-JUL-1998	40.475	-74.048	1			
R-EMAP Region 2 1998	1998	RB024	21-JUL-1998	40.475	-74.048	2	8.8	m	
R-EMAP Region 2 1993-94	1993	RB027	19-AUG-1993	40.471	-74.068	1	6.7	m	
R-EMAP Region 2 1998	1998	RB027	01-JUL-1998	40.471	-74.068	1			
R-EMAP Region 2 1998	1998	RB027	21-JUL-1998	40.471	-74.068	2	7.3	m	
R-EMAP Region 2 1993-94	1993	RB029	07-SEP-1993	40.465	-74.255	1	2.0	m	
R-EMAP Region 2 1998	1998	RB029	01-JUL-1998	40.464	-74.254	1			
R-EMAP Region 2 1998	1998	RB029	25-JUL-1998	40.464	-74.254	2	2.1	m	
R-EMAP Region 2 1993-94	1993	RB030	07-SEP-1993	40.455	-74.121	1	2.8	m	
R-EMAP Region 2 1998	1998	RB030	01-JUL-1998	40.455	-74.121	1			
R-EMAP Region 2 1998	1998	RB030	24-JUL-1998	40.455	-74.121	2	3.0	m	
R-EMAP Region 2 1993-94	1993	RB032	19-AUG-1993	40.447	-74.066	1	4.0	m	
R-EMAP Region 2 1998	1998	RB032	01-JUL-1998	40.447	-74.066	1			
R-EMAP Region 2 1998	1998	RB032	28-JUL-1998	40.447	-74.066	2	4.9	m	
R-EMAP Region 2 1993-94	1993	RB033	19-AUG-1993	40.438	-74.026	1	7.0	m	
R-EMAP Region 2 1998	1998	RB033	01-JUL-1998	40.439	-74.026	1			
R-EMAP Region 2 1998	1998	RB033	23-JUL-1998	40.439	-74.026	2	5.5	m	
R-EMAP Region 2 1993-94	1994	RB101	22-JUL-1994	40.587	-74.011	1	5.8	m	
R-EMAP Region 2 1993-94	1994	RB102	08-AUG-1994	40.573	-73.964	1	4.3	m	
R-EMAP Region 2 1993-94	1994	RB103	03-AUG-1994	40.558	-73.992	1	3.4	m	
R-EMAP Region 2 1993-94	1994	RB104	03-AUG-1994	40.55	-74.012	1	15.2	m	
R-EMAP Region 2 1993-94	1994	RB105	04-AUG-1994	40.541	-74.094	1	4.6	m	
R-EMAP Region 2 1993-94	1994	RB106	17-AUG-1994	40.514	-74.119	1	5.2	m	
R-EMAP Region 2 1993-94	1994	RB107	04-AUG-1994	40.513	-74.078	1	6.1	m	
R-EMAP Region 2 1993-94	1994	RB108	31-AUG-1994	40.513	-74.006	1	4.9	m	
R-EMAP Region 2 1993-94	1994	RB110	21-SEP-1994	40.486	-74.272	1	2.9	m	
R-EMAP Region 2 1993-94	1994	RB111	16-SEP-1994	40.475	-74.218	1	3.8	m	
R-EMAP Region 2 1993-94	1994	RB112	17-AUG-1994	40.472	-74.144	1	5.5	m	
R-EMAP Region 2 1993-94	1994	RB114	17-AUG-1994	40.468	-74.111	1	5.8	m	
R-EMAP Region 2 1993-94	1994	RB116	02-SEP-1994	40.486	-74.071	1	7.9	m	
R-EMAP Region 2 1993-94	1994	RB117	02-SEP-1994	40.464	-74.119	1	3.2	m	
R-EMAP Region 2 1998	1998	RB201	01-JUL-1998	40.574	-73.944	1			
R-EMAP Region 2 1998	1998	RB201	31-AUG-1998	40.574	-73.944	2	4.9	m	
R-EMAP Region 2 1998	1998	RB202	01-JUL-1998	40.515	-74.106	1			
R-EMAP Region 2 1998	1998	RB202	25-JUL-1998	40.515	-74.106	2	6.1	m	
R-EMAP Region 2 1998	1998	RB203	01-JUL-1998	40.426	-74.013	1			
R-EMAP Region 2 1998	1998	RB203	30-JUL-1998	40.426	-74.013	2	6.7	m	
R-EMAP Region 2 1998	1998	RB204	01-JUL-1998	40.48	-74.223	1			
R-EMAP Region 2 1998	1998	RB204	21-JUL-1998	40.48	-74.223	2			
R-EMAP Region 2 1998	1998	RB204	22-JUL-1998	40.48	-74.223	3	4.3	m	
R-EMAP Region 2 1998	1998	RB205	01-JUL-1998	40.455	-74.123	1			
R-EMAP Region 2 1998	1998	RB205	25-JUL-1998	40.455	-74.123	2	2.7	m	
R-EMAP Region 2 1998	1998	RB206	01-JUL-1998	40.544	-74.034	1			
R-EMAP Region 2 1998	1998	RB206	20-JUL-1998	40.544	-74.034	2	9.8	m	
R-EMAP Region 2 1998	1998	RB207	01-JUL-1998	40.587	-74.037	1			
R-EMAP Region 2 1998	1998	RB207	07-JUL-1998	40.587	-74.037	2	25.3	m	
R-EMAP Region 2 1998	1998	RB208	01-JUL-1998	40.498	-74.18	1			
R-EMAP Region 2 1998	1998	RB208	28-JUL-1998	40.498	-74.18	2	6.1	m	
R-EMAP Region 2 1998	1998	RB209	01-JUL-1998	40.516	-74.086	1			
R-EMAP Region 2 1998	1998	RB209	20-JUL-1998	40.516	-74.086	2	5.5	m	
R-EMAP Region 2 1998	1998	RB210	01-JUL-1998	40.477	-74.055	1			
R-EMAP Region 2 1998	1998	RB210	21-JUL-1998	40.477	-74.055	2	9.1	m	
R-EMAP Region 2 1998	1998	RB211	01-JUL-1998	40.461	-74.114	1			
R-EMAP Region 2 1998	1998	RB211	24-JUL-1998	40.461	-74.114	2	4.0	m	
R-EMAP Region 2 1998	1998	RB213	01-JUL-1998	40.585	-74.027	1			
R-EMAP Region 2 1998	1998	RB213	07-JUL-1998	40.585	-74.027	2	14.9	m	
R-EMAP Region 2 1998	1998	RB214	01-JUL-1998	40.547	-74.107	1			
R-EMAP Region 2 1998	1998	RB214	06-JUL-1998	40.547	-74.107	2	2.1	m	
R-EMAP Region 2 1998	1998	RB216	01-JUL-1998	40.471	-74.1	1			
R-EMAP Region 2 1998	1998	RB216	30-JUL-1998	40.471	-74.1	2	7.9	m	
R-EMAP Region 2 2003	2003	RB301	15-AUG-2003	40.588	-74.037	1	4.3	m	
R-EMAP Region 2 2003	2003	RB301	18-AUG-2003	40.588	-74.037	2	4.3	m	
R-EMAP Region 2 2003	2003	RB302	07-JUL-2003	40.586	-74.028	1	5.2	m	
R-EMAP Region 2 2003	2003	RB302	08-JUL-2003	40.586	-74.028	2	5.2	m	
R-EMAP Region 2 2003	2003	RB303	02-AUG-2003	40.582	-73.909	1	6.1	m	
R-EMAP Region 2 2003	2003	RB303	04-AUG-2003	40.582	-73.909	2	6.1	m	
R-EMAP Region 2 2003	2003	RB304	02-AUG-2003	40.575	-73.943	1	4.0	m	
R-EMAP Region 2 2003	2003	RB304	04-AUG-2003	40.575	-73.943	2	4.0	m	
R-EMAP Region 2 2003	2003	RB305	02-AUG-2003	40.498	-74.18	1	2.3	m	
R-EMAP Region 2 2003	2003	RB305	04-AUG-2003	40.498	-74.18	2	2.3	m	
R-EMAP Region 2 2003	2003	RB306	15-AUG-2003	40.546	-74.106	1	10.1	m	
R-EMAP Region 2 2003	2003	RB306	18-AUG-2003	40.546	-74.106	2	10.1	m	
R-EMAP Region 2 2003	2003	RB307	22-AUG-2003	40.528	-74.127	1	25.3	m	
R-EMAP Region 2 2003	2003	RB307	25-AUG-2003	40.528	-74.127	2	25.3	m	
R-EMAP Region 2 2003	2003	RB308	16-AUG-2003	40.515	-74.105	1	5.8	m	
R-EMAP Region 2 2003	2003	RB308	18-AUG-2003	40.515	-74.105	2	5.8	m	
R-EMAP Region 2 2003	2003	RB309	19-AUG-2003	40.516	-74.086	1	6.1	m	
R-EMAP Region 2 2003	2003	RB309	20-AUG-2003	40.516	-74.086	2	6.1	m	
R-EMAP Region 2 2003	2003	RB310	25-JUL-2003	40.513	-74.017	1	7.9	m	
R-EMAP Region 2 2003	2003	RB310	28-JUL-2003	40.513	-74.017	2	7.9	m	
R-EMAP Region 2 2003	2003	RB311	02-AUG-2003	40.431	-74.05	1	4.3	m	
R-EMAP Region 2 2003	2003	RB311	04-AUG-2003	40.431	-74.05	2	4.3	m	
R-EMAP Region 2 2003	2003	RB313	31-JUL-2003	40.426	-74.012	1	16.2	m	
R-EMAP Region 2 2003	2003	RB313	01-AUG-2003	40.426	-74.012	2	16.2	m	
R-EMAP Region 2 2003	2003	RB314	11-JUL-2003	40.477	-74.056	1	2.4	m	
R-EMAP Region 2 2003	2003	RB314	15-JUL-2003	40.477	-74.056	2	2.4	m	
R-EMAP Region 2 2003	2003	RB316	25-JUL-2003	40.478	-74.097	1	7.0	m	
R-EMAP Region 2 2003	2003	RB316	28-JUL-2003	40.478	-74.097	2	7.0	m	
R-EMAP Region 2 2003	2003	RB350	12-AUG-2003	40.457	-74.044	1	5.2	m	
R-EMAP Region 2 2003	2003	RB350	21-AUG-2003	40.457	-74.044	2	5.2	m	
R-EMAP Region 2 2003	2003	RB350	22-AUG-2003	40.457	-74.044	3	5.2	m	
R-EMAP Region 2 2003	2003	RB351	07-JUL-2003	40.481	-74.223	1	4.3	m	
R-EMAP Region 2 2003	2003	RB351	08-JUL-2003	40.481	-74.223	2	4.3	m	
R-EMAP Region 2 2003	2003	RB353	25-JUL-2003	40.46	-74.114	1	4.3	m	
R-EMAP Region 2 2003	2003	RB353	28-JUL-2003	40.46	-74.114	2	4.3	m	
R-EMAP Region 2 2003	2003	RB354	10-JUL-2003	40.477	-74.145	1	6.4	m	
R-EMAP Region 2 2003	2003	RB354	11-JUL-2003	40.477	-74.145	2	6.4	m	
R-EMAP Region 2 2003	2003	RB354	15-JUL-2003	40.477	-74.145	3	6.4	m	
R-EMAP Region 2 2003	2003	RB355	14-JUL-2003	40.472	-74.111	1	7.3	m	
R-EMAP Region 2 2003	2003	RB355	15-JUL-2003	40.472	-74.111	2	7.3	m	
R-EMAP Region 2 2003	2003	RB356	14-JUL-2003	40.455	-74.123	1	3.0	m	
R-EMAP Region 2 2003	2003	RB356	15-JUL-2003	40.455	-74.123	2	3.0	m	
R-EMAP Region 2 2003	2003	RB357	01-JUL-2003	40.557	-73.996	1	4.3	m	
R-EMAP Region 2 2003	2003	RB357	02-JUL-2003	40.557	-73.996	2	4.3	m	
R-EMAP Region 2 2003	2003	RB357	04-AUG-2003	40.557	-73.996	3	4.3	m	
R-EMAP Region 2 2003	2003	RB358	15-AUG-2003	40.512	-73.986	1	6.1	m	
R-EMAP Region 2 2003	2003	RB358	18-AUG-2003	40.512	-73.986	2	6.1	m	
R-EMAP Region 2 2003	2003	RB360	11-JUL-2003	40.526	-73.973	1	3.1	m	
R-EMAP Region 2 2003	2003	RB360	15-JUL-2003	40.526	-73.973	2	3.1	m	
R-EMAP Region 2 2003	2003	RB361	31-JUL-2003	40.545	-74.035	1	2.9	m	
R-EMAP Region 2 2003	2003	RB361	01-AUG-2003	40.545	-74.035	2	2.9	m	
R-EMAP Region 2 2003	2003	RB362	02-AUG-2003	40.516	-74.01	1	1.9	m	
R-EMAP Region 2 2003	2003	RB362	04-AUG-2003	40.516	-74.01	2	1.9	m	
R-EMAP Region 2 2003	2003	RB363	16-AUG-2003	40.511	-74.126	1	7.9	m	
R-EMAP Region 2 2003	2003	RB363	18-AUG-2003	40.511	-74.126	2	7.9	m	
R-EMAP Region 2 2003	2003	RB364	19-AUG-2003	40.445	-74.194	1	9.5	m	
R-EMAP Region 2 2003	2003	RB364	20-AUG-2003	40.445	-74.194	2	9.5	m	
R-EMAP Region 2 2003	2003	RB365	22-AUG-2003	40.425	-74.038	1	2.6	m	
R-EMAP Region 2 2003	2003	RB365	25-AUG-2003	40.425	-74.038	2	2.6	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0001-B	18-AUG-2000	41.466	-71.417	1	12.0	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0003-A	01-AUG-2000	41.479	-71.326	1	6.0	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0005-B	10-AUG-2000	41.508	-71.405	1	12.0	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0007-A	01-AUG-2000	41.494	-71.324	1	5.0	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0009-B	25-JUL-2000	41.473	-71.199	1	15.0	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0011-A	01-AUG-2000	41.515	-71.366	1	5.5	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0013-A	25-JUL-2000	41.514	-71.202	1	2.8	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0015-B	18-AUG-2000	41.567	-71.422	1	8.0	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0017-B	18-AUG-2000	41.554	-71.314	1	15.8	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0019-A	24-JUL-2000	41.559	-71.213	1	1.5	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0021-A	17-AUG-2000	41.597	-71.366	1	8.2	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0023-A	27-JUL-2000	41.596	-71.239	1	4.8	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0025-A	09-AUG-2000	41.659	-71.444	1	3.5	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0027-A	17-AUG-2000	41.621	-71.358	1	8.0	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0029-A	24-JUL-2000	41.614	-71.24	1	2.0	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0031-A	17-AUG-2000	41.667	-71.372	1	7.0	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0033-A	19-JUL-2000	41.666	-71.242	1	3.5	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0035-A	09-AUG-2000	41.696	-71.451	1	0.9	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0037-A	16-AUG-2000	41.708	-71.355	1	3.0	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0039-A	11-AUG-2000	41.701	-71.22	1	5.0	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0041-A	16-AUG-2000	41.73	-71.379	1	1.5	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0041-A	21-SEP-2000	41.73	-71.379	2	2.1	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0043-C	11-AUG-2000	41.722	-71.262	1	0.9	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0045-A	31-JUL-2000	41.771	-71.319	1	1.5	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0047-A	16-AUG-2000	41.825	-71.385	1	2.0	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0047-A	21-SEP-2000	41.825	-71.385	2	2.5	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0049-A	04-AUG-2000	41.318	-71.881	1	1.5	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0051-A	02-AUG-2000	41.332	-71.736	1	0.9	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0055-A	02-AUG-2000	41.379	-71.651	1	2.3	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0057-A	10-AUG-2000	41.381	-71.515	1	1.2	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0059-A	10-AUG-2000	41.4	-71.511	1	1.9	m	
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0061-A	08-AUG-2000	41.476	-71.381	2			
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0063-A	08-AUG-2000	41.462	-71.414	2			
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0065-A	11-AUG-2000	41.6	-71.23	2			
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0067-A	11-AUG-2000	41.68	-71.22	2			
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0069-A	10-AUG-2000	41.525	-71.342	2			
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0073-A	10-AUG-2000	41.551	-71.411	2			
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0075-A	09-AUG-2000	41.659	-71.375	2			
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0077-A	09-AUG-2000	41.67	-71.334	2			
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0081-A	10-AUG-2000	41.656	-71.238	2			
National Coastal Assessment-Northeast/Roger Williams University	2000	RI00-0083-A	11-AUG-2000	41.568	-71.219	2			
National Coastal Assessment-Northeast/University of Rhode Island	2001	RI01-0002-A	02-AUG-2001	41.471	-71.409	1	14.5	m	
National Coastal Assessment-Northeast/University of Rhode Island	2001	RI01-0004-B	01-AUG-2001	41.471	-71.206	1	14.5	m	
National Coastal Assessment-Northeast/University of Rhode Island	2001	RI01-0006-A	31-JUL-2001	41.507	-71.358	1	3.7	m	
National Coastal Assessment-Northeast/University of Rhode Island	2001	RI01-0008-A	01-AUG-2001	41.496	-71.222	1	10.9	m	
National Coastal Assessment-Northeast/University of Rhode Island	2001	RI01-0010-A	30-JUL-2001	41.54	-71.409	1	10.0	m	
National Coastal Assessment-Northeast/University of Rhode Island	2001	RI01-0012-A	31-JUL-2001	41.529	-71.319	1	12.2	m	
National Coastal Assessment-Northeast/University of Rhode Island	2001	RI01-0014-A	30-JUL-2001	41.578	-71.441	1	1.3	m	
National Coastal Assessment-Northeast/University of Rhode Island	2001	RI01-0016-A	20-JUL-2001	41.563	-71.359	1	10.6	m	
National Coastal Assessment-Northeast/University of Rhode Island	2001	RI01-0018-A	12-JUL-2001	41.566	-71.214	1	6.0	m	
National Coastal Assessment-Northeast/University of Rhode Island	2001	RI01-0020-A	30-JUL-2001	41.612	-71.407	1	8.5	m	
National Coastal Assessment-Northeast/University of Rhode Island	2001	RI01-0022-A	20-JUL-2001	41.61	-71.299	1	21.7	m	
National Coastal Assessment-Northeast/University of Rhode Island	2001	RI01-0024-A	12-JUL-2001	41.592	-71.21	1	3.6	m	
National Coastal Assessment-Northeast/University of Rhode Island	2001	RI01-0026-A	30-JUL-2001	41.641	-71.402	1	5.2	m	
National Coastal Assessment-Northeast/University of Rhode Island	2001	RI01-0028-A	12-JUL-2001	41.644	-71.272	1	7.6	m	
National Coastal Assessment-Northeast/University of Rhode Island	2001	RI01-0030-A	27-JUL-2001	41.667	-71.444	1	5.2	m	
National Coastal Assessment-Northeast/University of Rhode Island	2001	RI01-0032-A	16-JUL-2001	41.677	-71.339	1	7.5	m	
National Coastal Assessment-Northeast/University of Rhode Island	2001	RI01-0034-A	01-AUG-2001	41.683	-71.217	1	4.7	m	
National Coastal Assessment-Northeast/University of Rhode Island	2001	RI01-0036-A	27-JUL-2001	41.691	-71.39	1	1.4	m	
National Coastal Assessment-Northeast/University of Rhode Island	2001	RI01-0038-A	16-JUL-2001	41.701	-71.31	1	6.3	m	
National Coastal Assessment-Northeast/University of Rhode Island	2001	RI01-0040-A	11-JUL-2001	41.762	-71.318	1	1.5	m	
National Coastal Assessment-Northeast/University of Rhode Island	2001	RI01-0042-A	23-JUL-2001	41.801	-71.395	1	2.0	m	
National Coastal Assessment-Northeast/University of Rhode Island	2001	RI01-0044-B	11-JUL-2001	41.761	-71.285	1	2.5	m	
National Coastal Assessment-Northeast/University of Rhode Island	2001	RI01-0046-A	23-JUL-2001	41.81	-71.394	1	13.0	m	
National Coastal Assessment-Northeast/University of Rhode Island	2001	RI01-0048-A	23-JUL-2001	41.846	-71.372	1	2.2	m	
National Coastal Assessment-Northeast/University of Rhode Island	2001	RI01-0050-A	18-JUL-2001	41.318	-71.862	1	3.7	m	
National Coastal Assessment-Northeast/University of Rhode Island	2001	RI01-0052-A	17-JUL-2001	41.329	-71.786	1	0.4	m	
National Coastal Assessment-Northeast/University of Rhode Island	2001	RI01-0054-A	19-JUL-2001	41.367	-71.631	1	0.5	m	
National Coastal Assessment-Northeast/University of Rhode Island	2001	RI01-0056-A	19-JUL-2001	41.379	-71.645	1	1.5	m	
National Coastal Assessment-Northeast/University of Rhode Island	2001	RI01-0058-B	19-JUL-2001	41.396	-71.492	1	0.7	m	
National Coastal Assessment-Northeast/University of Rhode Island	2002	RI02-0056-B	25-SEP-2002	41.38	-71.647	1	4.1	m	
National Coastal Assessment-Northeast/University of Rhode Island	2002	RI02-0059-A	25-SEP-2002	41.4	-71.511	1	4.3	m	
National Coastal Assessment-Northeast/University of Rhode Island	2002	RI02-0061-A	18-JUL-2002	41.476	-71.381	1	3.7	m	
National Coastal Assessment-Northeast/University of Rhode Island	2002	RI02-0063-A	18-JUL-2002	41.462	-71.414	1	15.0	m	
National Coastal Assessment-Northeast/University of Rhode Island	2002	RI02-0065-A	16-JUL-2002	41.6	-71.23	1	5.5	m	
National Coastal Assessment-Northeast/University of Rhode Island	2002	RI02-0067-A	17-JUL-2002	41.68	-71.22	1	5.0	m	
National Coastal Assessment-Northeast/University of Rhode Island	2002	RI02-0069-A	17-JUL-2002	41.525	-71.342	1	8.5	m	
National Coastal Assessment-Northeast/University of Rhode Island	2002	RI02-0071-A	18-JUL-2002	41.596	-71.363	1	10.1	m	
National Coastal Assessment-Northeast/University of Rhode Island	2002	RI02-0073-A	19-JUL-2002	41.551	-71.411	1	2.4	m	
National Coastal Assessment-Northeast/University of Rhode Island	2002	RI02-0075-A	15-JUL-2002	41.659	-71.375	1	4.9	m	
National Coastal Assessment-Northeast/University of Rhode Island	2002	RI02-0077-A	15-JUL-2002	41.67	-71.334	1	1.8	m	
National Coastal Assessment-Northeast/University of Rhode Island	2002	RI02-0079-A	15-JUL-2002	41.705	-71.303	1	2.2	m	
National Coastal Assessment-Northeast/University of Rhode Island	2002	RI02-0081-A	17-JUL-2002	41.656	-71.238	1	6.7	m	
National Coastal Assessment-Northeast/University of Rhode Island	2002	RI02-0083-A	16-JUL-2002	41.568	-71.219	1	2.3	m	
National Coastal Assessment-Northeast/University of Rhode Island	2003	RI03-0301-A	26-AUG-2003	41.449	-71.373	1	26.6	m	
National Coastal Assessment-Northeast/University of Rhode Island	2003	RI03-0301-A	11-SEP-2003	41.449	-71.373	2	26.3	m	
National Coastal Assessment-Northeast/University of Rhode Island	2003	RI03-0302-A	14-AUG-2003	41.496	-71.414	1	12.5	m	
National Coastal Assessment-Northeast/University of Rhode Island	2003	RI03-0302-A	20-AUG-2003	41.496	-71.414	2	14.3	m	
National Coastal Assessment-Northeast/University of Rhode Island	2003	RI03-0306-A	28-JUL-2003	41.558	-71.408	1	7.8	m	
National Coastal Assessment-Northeast/University of Rhode Island	2003	RI03-0308-A	19-AUG-2003	41.561	-71.231	1	9.0	m	
National Coastal Assessment-Northeast/University of Rhode Island	2003	RI03-0311-A	27-AUG-2003	41.605	-71.291	1	21.4	m	
National Coastal Assessment-Northeast/University of Rhode Island	2003	RI03-0313-A	13-AUG-2003	41.626	-71.372	1	6.7	m	
National Coastal Assessment-Northeast/University of Rhode Island	2003	RI03-0316-A	07-AUG-2003	41.691	-71.348	1	6.1	m	
National Coastal Assessment-Northeast/University of Rhode Island	2003	RI03-0319-C	05-SEP-2003	41.812	-71.4	1	13.0	m	
National Coastal Assessment-Northeast/University of Rhode Island	2003	RI03-0321-A	20-AUG-2003	41.463	-71.388	1	6.6	m	
National Coastal Assessment-Northeast/University of Rhode Island	2003	RI03-0327-A	28-AUG-2003	41.579	-71.23	1	4.8	m	
National Coastal Assessment-Northeast/University of Rhode Island	2003	RI03-0329-A	06-AUG-2003	41.658	-71.39	1	3.5	m	
National Coastal Assessment-Northeast/University of Rhode Island	2003	RI03-0333-A	31-JUL-2003	41.72	-71.365	1	2.1	m	
National Coastal Assessment-Northeast/University of Rhode Island	2003	RI03-0334-A	12-AUG-2003	41.685	-71.217	1	1.7	m	
National Coastal Assessment-Northeast/University of Rhode Island	2003	RI03-0335-A	21-AUG-2003	41.703	-71.2	1	5.0	m	
National Coastal Assessment-Northeast/University of Rhode Island	2003	RI03-0337-C	05-SEP-2003	41.843	-71.372	1	2.5	m	
National Coastal Assessment-Northeast/University of Rhode Island	2003	RI03-0338-B	16-SEP-2003	41.325	-71.871	1	1.7	m	
National Coastal Assessment-Northeast/University of Rhode Island	2003	RI03-0361-A	16-JUL-2003	41.476	-71.381	1	10.1	m	
National Coastal Assessment-Northeast/University of Rhode Island	2003	RI03-0363-A	14-AUG-2003	41.462	-71.414	1	14.6	m	
National Coastal Assessment-Northeast/University of Rhode Island	2003	RI03-0367-A	15-JUL-2003	41.68	-71.22	1	5.1	m	
National Coastal Assessment-Northeast/University of Rhode Island	2003	RI03-0369-A	16-JUL-2003	41.525	-71.342	1	31.1	m	
National Coastal Assessment-Northeast/University of Rhode Island	2003	RI03-0371-A	14-JUL-2003	41.596	-71.363	1	6.7	m	
National Coastal Assessment-Northeast/University of Rhode Island	2003	RI03-0373-A	16-JUL-2003	41.551	-71.411	1	9.4	m	
National Coastal Assessment-Northeast/University of Rhode Island	2003	RI03-0375-A	07-AUG-2003	41.659	-71.375	1	19.2	m	
National Coastal Assessment-Northeast/University of Rhode Island	2003	RI03-0377-A	14-JUL-2003	41.67	-71.334	1	10.0	m	
National Coastal Assessment-Northeast/University of Rhode Island	2003	RI03-0379-A	14-JUL-2003	41.705	-71.303	1	5.5	m	
National Coastal Assessment-Northeast/University of Rhode Island	2003	RI03-0381-A	15-JUL-2003	41.656	-71.238	1	14.3	m	
National Coastal Assessment-Northeast/University of Rhode Island	2003	RI03-0383-A	15-JUL-2003	41.568	-71.219	1	8.5	m	
National Coastal Assessment-Northeast/University of Rhode Island	2004	RI04-0304-A	22-JUL-2004	41.498	-71.325	1	7.2	m	
National Coastal Assessment-Northeast/University of Rhode Island	2004	RI04-0307-A	09-AUG-2004	41.566	-71.344	1	10.0	m	
National Coastal Assessment-Northeast/University of Rhode Island	2004	RI04-0314-A	03-AUG-2004	41.641	-71.3	1	11.0	m	
National Coastal Assessment-Northeast/University of Rhode Island	2004	RI04-0317-A	03-AUG-2004	41.7	-71.314	1	7.2	m	
National Coastal Assessment-Northeast/University of Rhode Island	2004	RI04-0320-B	29-JUL-2004	41.817	-71.393	1	5.8	m	
National Coastal Assessment-Northeast/University of Rhode Island	2004	RI04-0322-A	02-AUG-2004	41.467	-71.429	1	5.0	m	
National Coastal Assessment-Northeast/University of Rhode Island	2004	RI04-0324-B	21-JUL-2004	41.488	-71.243	1	3.0	m	
National Coastal Assessment-Northeast/University of Rhode Island	2004	RI04-0326-A	08-JUL-2004	41.572	-71.431	1	4.2	m	
National Coastal Assessment-Northeast/University of Rhode Island	2004	RI04-0328-A	21-JUL-2004	41.578	-71.209	1	2.0	m	
National Coastal Assessment-Northeast/University of Rhode Island	2004	RI04-0329-A	12-JUL-2004	41.658	-71.39	1	3.6	m	
National Coastal Assessment-Northeast/University of Rhode Island	2004	RI04-0330-A	06-JUL-2004	41.647	-71.37	1	7.1	m	
National Coastal Assessment-Northeast/University of Rhode Island	2004	RI04-0330-A	09-JUL-2004	41.647	-71.37	2	7.0	m	
National Coastal Assessment-Northeast/University of Rhode Island	2004	RI04-0332-A	09-JUL-2004	41.685	-71.448	1	2.4	m	
National Coastal Assessment-Northeast/University of Rhode Island	2004	RI04-0333-A	02-JUL-2004	41.72	-71.365	1	2.7	m	
National Coastal Assessment-Northeast/University of Rhode Island	2004	RI04-0333-A	09-JUL-2004	41.72	-71.365	2	1.9	m	
National Coastal Assessment-Northeast/University of Rhode Island	2004	RI04-0335-A	19-JUL-2004	41.703	-71.2	1	5.6	m	
National Coastal Assessment-Northeast/University of Rhode Island	2004	RI04-0336-A	30-JUL-2004	41.76	-71.305	1	0.9	m	
National Coastal Assessment-Northeast/University of Rhode Island	2004	RI04-0339-A	12-AUG-2004	41.356	-71.671	1	1.2	m	
National Coastal Assessment-Northeast/University of Rhode Island	2004	RI04-0461-A	21-JUL-2004	41.476	-71.381	1	11.5	m	
National Coastal Assessment-Northeast/University of Rhode Island	2004	RI04-0463-A	19-JUL-2004	41.462	-71.414	1	13.9	m	
National Coastal Assessment-Northeast/University of Rhode Island	2004	RI04-0467-A	20-JUL-2004	41.68	-71.22	1	5.8	m	
National Coastal Assessment-Northeast/University of Rhode Island	2004	RI04-0469-A	16-JUL-2004	41.525	-71.342	1	29.7	m	
National Coastal Assessment-Northeast/University of Rhode Island	2004	RI04-0471-A	11-AUG-2004	41.596	-71.363	1	7.0	m	
National Coastal Assessment-Northeast/University of Rhode Island	2004	RI04-0473-A	11-AUG-2004	41.551	-71.411	1	11.0	m	
National Coastal Assessment-Northeast/University of Rhode Island	2004	RI04-0475-A	14-JUL-2004	41.659	-71.375	1	21.3	m	
National Coastal Assessment-Northeast/University of Rhode Island	2004	RI04-0477-A	14-JUL-2004	41.67	-71.334	1	6.1	m	
National Coastal Assessment-Northeast/University of Rhode Island	2004	RI04-0481-A	20-JUL-2004	41.656	-71.238	1	15.2	m	
National Coastal Assessment-Northeast/University of Rhode Island	2004	RI04-0483-A	20-JUL-2004	41.568	-71.219	1	9.8	m	
National Coastal Assessment-Northeast/University of Rhode Island	2004	RI04-0486-A	21-JUL-2004	41.461	-71.377	1	31.7	m	
National Coastal Assessment-Northeast/University of Rhode Island	2004	RI04-0487-A	20-JUL-2004	41.501	-71.216	1	8.5	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0001-A	15-AUG-2005	41.604	-71.294	1	22.4	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0002-A	01-AUG-2005	41.606	-71.235	1	4.2	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0003-A	05-JUL-2005	41.703	-71.2	1	4.7	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0004-C	18-AUG-2005	41.525	-71.326	1	16.0	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0005-A	28-JUL-2005	41.622	-71.413	1	4.4	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0006-C	09-AUG-2005	41.483	-71.341	1	23.5	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0007-A	10-AUG-2005	41.655	-71.307	1	11.4	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0008-A	01-AUG-2005	41.484	-71.228	1	13.3	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0009-A	01-JUL-2005	41.52	-71.224	1	6.2	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0010-A	06-JUL-2005	41.519	-71.363	1	1.6	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0011-A	19-JUL-2005	41.687	-71.298	1	4.2	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0012-A	19-JUL-2005	41.62	-71.36	1	7.8	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0013-A	12-JUL-2005	41.658	-71.39	1	4.4	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0014-A	03-AUG-2005	41.478	-71.363	1	6.4	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0015-A	21-JUL-2005	41.627	-71.286	1	11.8	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0016-A	16-AUG-2005	41.328	-71.79	1	0.4	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0017-A	27-JUL-2005	41.801	-71.393	1	1.9	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0018-A	29-JUL-2005	41.387	-71.513	1	1.0	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0018-A	24-AUG-2005	41.387	-71.513	2	2.8	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0019-A	13-JUL-2005	41.72	-71.365	1	2.8	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0019-A	10-AUG-2005	41.72	-71.365	2	3.4	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0020-A	05-AUG-2005	41.452	-71.411	1	17.9	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0021-A	15-JUL-2005	41.636	-71.269	1	9.4	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0022-A	08-AUG-2005	41.54	-71.352	1	20.3	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0023-A	26-JUL-2005	41.719	-71.29	1	1.9	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0024-A	18-JUL-2005	41.578	-71.341	1	9.8	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0025-A	05-JUL-2005	41.709	-71.165	1	7.0	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0561-A	12-JUL-2005	41.476	-71.381	1	11.2	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0563-A	15-JUL-2005	41.462	-71.414	1	13.1	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0567-A	13-JUL-2005	41.68	-71.22	1	4.9	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0567-A	18-AUG-2005	41.68	-71.22	2	3.6	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0569-A	15-JUL-2005	41.525	-71.342	1	22.0	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0571-A	11-JUL-2005	41.596	-71.363	1	8.0	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0573-A	15-JUL-2005	41.551	-71.411	1	9.8	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0575-A	19-AUG-2005	41.659	-71.375	1	16.1	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0577-A	11-JUL-2005	41.67	-71.334	1	6.7	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0581-A	13-JUL-2005	41.656	-71.238	1	11.0	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0583-A	13-JUL-2005	41.568	-71.219	1	10.4	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0586-A	19-AUG-2005	41.461	-71.377	1	25.9	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0587-A	13-JUL-2005	41.501	-71.216	1	8.8	m	
National Coastal Assessment-Northeast/University of Rhode Island	2005	RI05-0587-A	18-AUG-2005	41.501	-71.216	2	9.2	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0026-A	11-AUG-2006	41.846	-71.37	1	2.0	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0027-B	05-JUL-2006	41.643	-71.343	1	2.0	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0027-B	06-JUL-2006	41.643	-71.343	2	1.1	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0028-A	08-AUG-2006	41.72	-71.365	1	3.0	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0029-A	19-JUL-2006	41.463	-71.413	1	13.4	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0030-A	25-JUL-2006	41.658	-71.253	1	4.3	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0030-A	31-JUL-2006	41.658	-71.253	2	4.5	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0031-A	11-JUL-2006	41.577	-71.421	1	4.5	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0031-A	12-JUL-2006	41.577	-71.421	2	5.5	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0032-A	31-JUL-2006	41.698	-71.324	1	8.0	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0033-A	11-JUL-2006	41.611	-71.41	1	2.4	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0034-B	11-AUG-2006	41.76	-71.308	1	1.4	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0035-A	07-AUG-2006	41.367	-71.645	1	1.4	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0036-A	15-AUG-2006	41.625	-71.337	1	6.1	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0037-A	17-JUL-2006	41.469	-71.228	1	17.7	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0037-A	09-AUG-2006	41.469	-71.228	2	18.0	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0038-A	07-JUL-2006	41.631	-71.234	1	0.8	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0038-A	10-JUL-2006	41.631	-71.234	2	0.8	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0039-A	24-JUL-2006	41.546	-71.32	1	16.7	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0040-A	07-JUL-2006	41.575	-71.227	1	4.6	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0041-A	26-JUL-2006	41.578	-71.379	1	8.5	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0042-A	02-AUG-2006	41.58	-71.307	1	16.8	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0042-A	09-AUG-2006	41.58	-71.307	2	18.3	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0043-A	14-AUG-2006	41.555	-71.393	1	9.8	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0044-A	10-JUL-2006	41.703	-71.2	1	5.0	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0045-A	25-JUL-2006	41.528	-71.345	1	9.5	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0046-A	16-AUG-2006	41.658	-71.39	1	3.7	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0047-A	26-JUL-2006	41.508	-71.385	1	3.6	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0048-A	06-JUL-2006	41.621	-71.305	1	1.6	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0049-A	03-AUG-2006	41.478	-71.201	1	12.0	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0050-A	18-JUL-2006	41.538	-71.235	1	1.4	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0661-A	12-JUL-2006	41.476	-71.381	1	13.4	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0663-A	12-JUL-2006	41.462	-71.414	1	15.1	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0667-A	11-JUL-2006	41.68	-71.22	1	4.5	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0669-A	10-JUL-2006	41.525	-71.342	1	22.9	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0671-A	10-JUL-2006	41.596	-71.363	1	7.8	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0671-A	17-AUG-2006	41.596	-71.363	2	6.9	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0673-A	17-AUG-2006	41.551	-71.411	1	9.1	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0675-A	10-JUL-2006	41.659	-71.375	1	21.3	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0675-A	17-AUG-2006	41.659	-71.375	2	23.6	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0677-A	10-JUL-2006	41.67	-71.334	1	6.2	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0677-A	17-AUG-2006	41.67	-71.334	2	5.9	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0681-A	11-JUL-2006	41.656	-71.238	1	14.0	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0683-A	11-JUL-2006	41.568	-71.219	1	7.4	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0686-A	12-JUL-2006	41.461	-71.377	1	36.7	m	
National Coastal Assessment-Northeast/University of Rhode Island	2006	RI06-0687-A	11-JUL-2006	41.501	-71.216	1	10.0	m	
DE/MD Coastal Bays	1993	STN_1	01-JUL-1993	38.596	-75.288	1			
DE/MD Coastal Bays	1993	STN_1	01-AUG-1993	38.596	-75.288	2			
DE/MD Coastal Bays	1993	STN_1	01-SEP-1993	38.596	-75.288	3			
DE/MD Coastal Bays	1993	STN_10	01-JUL-1993	38.593	-75.197	1			
DE/MD Coastal Bays	1993	STN_10	01-AUG-1993	38.593	-75.197	2			
DE/MD Coastal Bays	1993	STN_10	01-SEP-1993	38.593	-75.197	3			
DE/MD Coastal Bays	1993	STN_11	01-JUL-1993	38.579	-75.184	1			
DE/MD Coastal Bays	1993	STN_11	01-AUG-1993	38.579	-75.184	2			
DE/MD Coastal Bays	1993	STN_11	01-SEP-1993	38.579	-75.184	3			
DE/MD Coastal Bays	1993	STN_12	01-JUL-1993	38.583	-75.182	1			
DE/MD Coastal Bays	1993	STN_12	01-AUG-1993	38.583	-75.182	2			
DE/MD Coastal Bays	1993	STN_12	01-SEP-1993	38.583	-75.182	3			
DE/MD Coastal Bays	1993	STN_13	01-JUL-1993	38.576	-75.185	1			
DE/MD Coastal Bays	1993	STN_13	01-AUG-1993	38.576	-75.185	2			
DE/MD Coastal Bays	1993	STN_13	01-SEP-1993	38.576	-75.185	3			
DE/MD Coastal Bays	1993	STN_14	01-JUL-1993	38.603	-75.157	1			
DE/MD Coastal Bays	1993	STN_14	01-AUG-1993	38.603	-75.157	2			
DE/MD Coastal Bays	1993	STN_14	01-SEP-1993	38.603	-75.157	3			
DE/MD Coastal Bays	1993	STN_15	01-JUL-1993	38.588	-75.153	1			
DE/MD Coastal Bays	1993	STN_15	01-AUG-1993	38.588	-75.153	2			
DE/MD Coastal Bays	1993	STN_15	01-SEP-1993	38.588	-75.153	3			
DE/MD Coastal Bays	1993	STN_16	01-JUL-1993	38.576	-75.099	1			
DE/MD Coastal Bays	1993	STN_16	01-AUG-1993	38.576	-75.099	2			
DE/MD Coastal Bays	1993	STN_16	01-SEP-1993	38.576	-75.099	3			
DE/MD Coastal Bays	1993	STN_18	01-JUL-1993	38.603	-75.079	1			
DE/MD Coastal Bays	1993	STN_18	01-AUG-1993	38.603	-75.079	2			
DE/MD Coastal Bays	1993	STN_18	01-SEP-1993	38.603	-75.079	3			
DE/MD Coastal Bays	1993	STN_19	01-JUL-1993	38.611	-75.086	1			
DE/MD Coastal Bays	1993	STN_19	01-AUG-1993	38.611	-75.086	2			
DE/MD Coastal Bays	1993	STN_19	01-SEP-1993	38.611	-75.086	3			
DE/MD Coastal Bays	1993	STN_2	01-JUL-1993	38.59	-75.27	1			
DE/MD Coastal Bays	1993	STN_2	01-AUG-1993	38.59	-75.27	2			
DE/MD Coastal Bays	1993	STN_2	01-SEP-1993	38.59	-75.27	3			
DE/MD Coastal Bays	1993	STN_20	01-JUL-1993	38.618	-75.101	1			
DE/MD Coastal Bays	1993	STN_20	01-AUG-1993	38.618	-75.101	2			
DE/MD Coastal Bays	1993	STN_20	01-SEP-1993	38.618	-75.101	3			
DE/MD Coastal Bays	1993	STN_21	01-JUL-1993	38.615	-75.121	1			
DE/MD Coastal Bays	1993	STN_21	01-AUG-1993	38.615	-75.121	2			
DE/MD Coastal Bays	1993	STN_21	01-SEP-1993	38.615	-75.121	3			
DE/MD Coastal Bays	1993	STN_22	01-JUL-1993	38.634	-75.109	1			
DE/MD Coastal Bays	1993	STN_22	01-AUG-1993	38.634	-75.109	2			
DE/MD Coastal Bays	1993	STN_22	01-SEP-1993	38.634	-75.109	3			
DE/MD Coastal Bays	1993	STN_23	01-JUL-1993	38.639	-75.082	1			
DE/MD Coastal Bays	1993	STN_24	01-JUL-1993	38.635	-75.125	1			
DE/MD Coastal Bays	1993	STN_24	01-AUG-1993	38.635	-75.125	2			
DE/MD Coastal Bays	1993	STN_24	01-SEP-1993	38.635	-75.125	3			
DE/MD Coastal Bays	1993	STN_25	01-JUL-1993	38.654	-75.127	1			
DE/MD Coastal Bays	1993	STN_25	01-AUG-1993	38.654	-75.127	2			
DE/MD Coastal Bays	1993	STN_25	01-SEP-1993	38.654	-75.127	3			
DE/MD Coastal Bays	1993	STN_26	01-JUL-1993	38.688	-75.133	1			
DE/MD Coastal Bays	1993	STN_26	01-AUG-1993	38.688	-75.133	2			
DE/MD Coastal Bays	1993	STN_26	01-SEP-1993	38.688	-75.133	3			
DE/MD Coastal Bays	1993	STN_27	01-JUL-1993	38.691	-75.1	1			
DE/MD Coastal Bays	1993	STN_27	01-AUG-1993	38.691	-75.1	2			
DE/MD Coastal Bays	1993	STN_27	01-SEP-1993	38.691	-75.1	3			
DE/MD Coastal Bays	1993	STN_28	01-JUL-1993	38.687	-75.076	1			
DE/MD Coastal Bays	1993	STN_28	01-AUG-1993	38.687	-75.076	2			
DE/MD Coastal Bays	1993	STN_28	01-SEP-1993	38.687	-75.076	3			
DE/MD Coastal Bays	1993	STN_29	01-JUL-1993	38.687	-75.076	1			
DE/MD Coastal Bays	1993	STN_29	01-AUG-1993	38.687	-75.076	2			
DE/MD Coastal Bays	1993	STN_29	01-SEP-1993	38.687	-75.076	3			
DE/MD Coastal Bays	1993	STN_3	01-JUL-1993	38.59	-75.25	1			
DE/MD Coastal Bays	1993	STN_3	01-AUG-1993	38.59	-75.25	2			
DE/MD Coastal Bays	1993	STN_3	01-SEP-1993	38.59	-75.25	3			
DE/MD Coastal Bays	1993	STN_4	01-JUL-1993	38.593	-75.247	1			
DE/MD Coastal Bays	1993	STN_4	01-AUG-1993	38.593	-75.247	2			
DE/MD Coastal Bays	1993	STN_4	01-SEP-1993	38.593	-75.247	3			
DE/MD Coastal Bays	1993	STN_5	01-JUL-1993	38.588	-75.227	1			
DE/MD Coastal Bays	1993	STN_5	01-AUG-1993	38.588	-75.227	2			
DE/MD Coastal Bays	1993	STN_5	01-SEP-1993	38.588	-75.227	3			
DE/MD Coastal Bays	1993	STN_6	01-JUL-1993	38.591	-75.226	1			
DE/MD Coastal Bays	1993	STN_6	01-AUG-1993	38.591	-75.226	2			
DE/MD Coastal Bays	1993	STN_6	01-SEP-1993	38.591	-75.226	3			
DE/MD Coastal Bays	1993	STN_7	01-JUL-1993	38.591	-75.213	1			
DE/MD Coastal Bays	1993	STN_7	01-AUG-1993	38.591	-75.213	2			
DE/MD Coastal Bays	1993	STN_7	01-SEP-1993	38.591	-75.213	3			
DE/MD Coastal Bays	1993	STN_9	01-JUL-1993	38.586	-75.205	1			
DE/MD Coastal Bays	1993	STN_9	01-AUG-1993	38.586	-75.205	2			
DE/MD Coastal Bays	1993	STN_9	01-SEP-1993	38.586	-75.205	3			
R-EMAP Region 2 1993-94	1993	UH003	24-AUG-1993	40.868	-73.944	1	8.5	m	
R-EMAP Region 2 1998	1998	UH003	01-JUN-1998	40.867	-73.944	1			
R-EMAP Region 2 1998	1998	UH003	01-JUL-1998	40.867	-73.944	2	9.1	m	
R-EMAP Region 2 1993-94	1993	UH004	24-AUG-1993	40.865	-73.941	1	12.5	m	
R-EMAP Region 2 1998	1998	UH004	01-JUN-1998	40.865	-73.94	1			
R-EMAP Region 2 1998	1998	UH004	01-JUL-1998	40.865	-73.94	2	13.4	m	
R-EMAP Region 2 1993-94	1993	UH008	31-AUG-1993	40.802	-73.813	1	14.6	m	
R-EMAP Region 2 1998	1998	UH008	01-JUN-1998	40.802	-73.813	1			
R-EMAP Region 2 1998	1998	UH008	24-AUG-1998	40.802	-73.813	2	13.7	m	
R-EMAP Region 2 1993-94	1993	UH010	31-AUG-1993	40.791	-73.896	1	4.9	m	
R-EMAP Region 2 1998	1998	UH010	01-JUN-1998	40.791	-73.897	1			
R-EMAP Region 2 1998	1998	UH010	26-AUG-1998	40.791	-73.897	2	6.7	m	
R-EMAP Region 2 1993-94	1993	UH011	10-SEP-1993	40.785	-73.874	1	2.6	m	
R-EMAP Region 2 1998	1998	UH011	01-JUN-1998	40.786	-73.874	1			
R-EMAP Region 2 1998	1998	UH011	09-JUL-1998	40.786	-73.874	2	3.0	m	
R-EMAP Region 2 1993-94	1993	UH014	25-AUG-1993	40.756	-74.02	1	7.6	m	
R-EMAP Region 2 1998	1998	UH014	01-JUN-1998	40.756	-74.02	1			
R-EMAP Region 2 1998	1998	UH014	22-AUG-1998	40.756	-74.02	2	7.0	m	
R-EMAP Region 2 1993-94	1993	UH018	25-AUG-1993	40.707	-74.022	1	17.1	m	
R-EMAP Region 2 1998	1998	UH018	01-JUN-1998	40.707	-74.022	1			
R-EMAP Region 2 1998	1998	UH018	03-JUL-1998	40.707	-74.022	2	14.6	m	
R-EMAP Region 2 1993-94	1993	UH019	21-SEP-1993	40.691	-74.041	1	7.6	m	
R-EMAP Region 2 1998	1998	UH019	01-JUN-1998	40.691	-74.04	1			
R-EMAP Region 2 1998	1998	UH019	03-JUL-1998	40.691	-74.04	2	8.8	m	
R-EMAP Region 2 1993-94	1993	UH020	26-AUG-1993	40.689	-74.004	1	11.6	m	
R-EMAP Region 2 1998	1998	UH020	01-JUN-1998	40.69	-74.004	1			
R-EMAP Region 2 1998	1998	UH020	28-AUG-1998	40.69	-74.004	2	11.0	m	
R-EMAP Region 2 1993-94	1993	UH022	03-SEP-1993	40.677	-74.047	1	9.1	m	
R-EMAP Region 2 1998	1998	UH022	01-JUN-1998	40.676	-74.046	1			
R-EMAP Region 2 1998	1998	UH022	23-JUN-1998	40.676	-74.046	2	15.8	m	
R-EMAP Region 2 1993-94	1993	UH023	02-SEP-1993	40.663	-74.029	1	4.6	m	
R-EMAP Region 2 1998	1998	UH023	01-JUN-1998	40.664	-74.028	1			
R-EMAP Region 2 1998	1998	UH023	23-JUN-1998	40.664	-74.028	2	4.6	m	
R-EMAP Region 2 1993-94	1993	UH026	21-SEP-1993	40.654	-74.043	1	12.5	m	
R-EMAP Region 2 1998	1998	UH026	01-JUN-1998	40.655	-74.043	1			
R-EMAP Region 2 1998	1998	UH026	26-JUN-1998	40.655	-74.043	2	12.5	m	
R-EMAP Region 2 1993-94	1993	UH029	20-AUG-1993	40.636	-74.052	1	14.6	m	
R-EMAP Region 2 1998	1998	UH029	01-JUN-1998	40.636	-74.051	1			
R-EMAP Region 2 1998	1998	UH029	27-JUN-1998	40.636	-74.051	2	4.6	m	
R-EMAP Region 2 1993-94	1993	UH030	20-AUG-1993	40.62	-74.06	1	24.4	m	
R-EMAP Region 2 1998	1998	UH030	01-JUN-1998	40.619	-74.06	1			
R-EMAP Region 2 1998	1998	UH030	02-JUL-1998	40.619	-74.06	2	23.8	m	
R-EMAP Region 2 1993-94	1994	UH101	14-AUG-1994	40.687	-74.027	1	15.2	m	
R-EMAP Region 2 1993-94	1994	UH102	14-AUG-1994	40.914	-73.923	1	7.9	m	
R-EMAP Region 2 1993-94	1994	UH103	14-AUG-1994	40.891	-73.934	1	5.5	m	
R-EMAP Region 2 1993-94	1994	UH104	01-SEP-1994	40.811	-73.814	1	4.0	m	
R-EMAP Region 2 1993-94	1994	UH105	14-AUG-1994	40.803	-73.98	1	16.5	m	
R-EMAP Region 2 1993-94	1994	UH106	13-AUG-1994	40.796	-73.875	1	13.7	m	
R-EMAP Region 2 1993-94	1994	UH107	01-SEP-1994	40.796	-73.895	1	9.1	m	
R-EMAP Region 2 1993-94	1994	UH108	14-AUG-1994	40.714	-74.029	1	11.6	m	
R-EMAP Region 2 1993-94	1994	UH109	19-AUG-1994	40.696	-74.064	1	3.4	m	
R-EMAP Region 2 1993-94	1994	UH110	27-JUL-1994	40.681	-74.05	1	2.3	m	
R-EMAP Region 2 1993-94	1994	UH111	13-AUG-1994	40.68	-74.041	1	18.9	m	
R-EMAP Region 2 1993-94	1994	UH112	19-AUG-1994	40.674	-74.091	1	3.4	m	
R-EMAP Region 2 1993-94	1994	UH113	27-JUL-1994	40.658	-74.077	1	3.9	m	
R-EMAP Region 2 1993-94	1994	UH114	13-AUG-1994	40.649	-74.055	1	15.5	m	
R-EMAP Region 2 1998	1998	UH201	01-JUN-1998	40.665	-74.013	1			
R-EMAP Region 2 1998	1998	UH201	25-AUG-1998	40.665	-74.013	2	11.6	m	
R-EMAP Region 2 1998	1998	UH202	01-JUN-1998	40.616	-74.061	1			
R-EMAP Region 2 1998	1998	UH202	24-JUN-1998	40.616	-74.061	2	19.2	m	
R-EMAP Region 2 1998	1998	UH204	01-JUN-1998	40.864	-73.939	1			
R-EMAP Region 2 1998	1998	UH204	03-JUL-1998	40.864	-73.939	2	14.3	m	
R-EMAP Region 2 1998	1998	UH206	01-JUN-1998	40.776	-73.888	1			
R-EMAP Region 2 1998	1998	UH206	09-JUL-1998	40.776	-73.888	2	4.3	m	
R-EMAP Region 2 1998	1998	UH208	01-JUN-1998	40.676	-74.042	1			
R-EMAP Region 2 1998	1998	UH208	26-JUN-1998	40.676	-74.042	2	19.2	m	
R-EMAP Region 2 1998	1998	UH209	01-JUN-1998	40.623	-74.066	1			
R-EMAP Region 2 1998	1998	UH209	27-JUN-1998	40.623	-74.066	2	4.0	m	
R-EMAP Region 2 1998	1998	UH211	01-JUN-1998	40.851	-73.951	1			
R-EMAP Region 2 1998	1998	UH211	29-JUN-1998	40.851	-73.951	2	4.9	m	
R-EMAP Region 2 1998	1998	UH212	01-JUN-1998	40.803	-73.811	1			
R-EMAP Region 2 1998	1998	UH212	24-AUG-1998	40.803	-73.811	2	16.2	m	
R-EMAP Region 2 1998	1998	UH213	01-JUN-1998	40.773	-73.999	1			
R-EMAP Region 2 1998	1998	UH213	22-AUG-1998	40.773	-73.999	2	13.4	m	
R-EMAP Region 2 1998	1998	UH214	01-JUN-1998	40.681	-74.061	1			
R-EMAP Region 2 1998	1998	UH214	22-JUN-1998	40.681	-74.061	2	2.6	m	
R-EMAP Region 2 1998	1998	UH215	01-JUN-1998	40.638	-74.064	1			
R-EMAP Region 2 1998	1998	UH215	12-AUG-1998	40.638	-74.064	2	17.1	m	
R-EMAP Region 2 1998	1998	UH216	01-JUN-1998	40.712	-74.024	1			
R-EMAP Region 2 1998	1998	UH216	12-AUG-1998	40.712	-74.024	2	17.1	m	
R-EMAP Region 2 1998	1998	UH217	01-JUN-1998	40.808	-73.828	1			
R-EMAP Region 2 1998	1998	UH217	27-AUG-1998	40.808	-73.828	2	2.1	m	
R-EMAP Region 2 1998	1998	UH219	01-JUN-1998	40.695	-74.037	1			
R-EMAP Region 2 1998	1998	UH219	28-AUG-1998	40.695	-74.037	2	8.5	m	
R-EMAP Region 2 2003	2003	UH301	09-JUL-2003	40.785	-73.993	1	7.0	m	
R-EMAP Region 2 2003	2003	UH302	22-JUL-2003	40.773	-73.998	1	16.2	m	
R-EMAP Region 2 2003	2003	UH302	23-JUL-2003	40.773	-73.998	2	16.2	m	
R-EMAP Region 2 2003	2003	UH304	28-AUG-2003	40.695	-74.037	1	15.5	m	
R-EMAP Region 2 2003	2003	UH304	29-AUG-2003	40.695	-74.037	2	15.5	m	
R-EMAP Region 2 2003	2003	UH308	23-AUG-2003	40.665	-74.013	1	17.4	m	
R-EMAP Region 2 2003	2003	UH308	25-AUG-2003	40.665	-74.013	2	17.4	m	
R-EMAP Region 2 2003	2003	UH309	22-JUL-2003	40.675	-74.044	1	15.5	m	
R-EMAP Region 2 2003	2003	UH309	24-JUL-2003	40.675	-74.044	2	15.5	m	
R-EMAP Region 2 2003	2003	UH309	25-JUL-2003	40.675	-74.044	3	15.5	m	
R-EMAP Region 2 2003	2003	UH311	20-AUG-2003	40.681	-74.06	1	13.7	m	
R-EMAP Region 2 2003	2003	UH311	21-AUG-2003	40.681	-74.06	2	13.7	m	
R-EMAP Region 2 2003	2003	UH312	01-AUG-2003	40.659	-74.065	1	12.5	m	
R-EMAP Region 2 2003	2003	UH312	04-AUG-2003	40.659	-74.065	2	12.5	m	
R-EMAP Region 2 2003	2003	UH313	25-AUG-2003	40.616	-74.061	1	9.8	m	
R-EMAP Region 2 2003	2003	UH313	28-AUG-2003	40.616	-74.061	2	9.8	m	
R-EMAP Region 2 2003	2003	UH313	29-AUG-2003	40.616	-74.061	3	9.8	m	
R-EMAP Region 2 2003	2003	UH314	24-JUL-2003	40.623	-74.065	1	2.6	m	
R-EMAP Region 2 2003	2003	UH314	25-JUL-2003	40.623	-74.065	2	2.6	m	
R-EMAP Region 2 2003	2003	UH315	23-AUG-2003	40.639	-74.064	1	16.5	m	
R-EMAP Region 2 2003	2003	UH315	25-AUG-2003	40.639	-74.064	2	16.5	m	
R-EMAP Region 2 2003	2003	UH316	23-AUG-2003	40.649	-74.037	1	15.9	m	
R-EMAP Region 2 2003	2003	UH316	25-AUG-2003	40.649	-74.037	2	15.9	m	
R-EMAP Region 2 2003	2003	UH319	24-JUL-2003	40.736	-73.967	1	6.7	m	
R-EMAP Region 2 2003	2003	UH319	25-JUL-2003	40.736	-73.967	2	6.7	m	
R-EMAP Region 2 2003	2003	UH351	04-AUG-2003	40.757	-73.959	1	12.5	m	
R-EMAP Region 2 2003	2003	UH351	05-AUG-2003	40.757	-73.959	2	12.5	m	
R-EMAP Region 2 2003	2003	UH352	23-AUG-2003	40.711	-74.024	1	15.5	m	
R-EMAP Region 2 2003	2003	UH352	25-AUG-2003	40.711	-74.024	2	15.5	m	
R-EMAP Region 2 2003	2003	UH352	29-AUG-2003	40.711	-74.024	3	15.5	m	
R-EMAP Region 2 2003	2003	UH354	21-JUL-2003	40.905	-73.929	1	12.8	m	
R-EMAP Region 2 2003	2003	UH355	20-AUG-2003	40.864	-73.94	1	16.2	m	
R-EMAP Region 2 2003	2003	UH355	21-AUG-2003	40.864	-73.94	2	16.2	m	
R-EMAP Region 2 2003	2003	UH356	25-AUG-2003	40.85	-73.951	1	2.7	m	
R-EMAP Region 2 2003	2003	UH356	26-AUG-2003	40.85	-73.951	2	2.7	m	
R-EMAP Region 2 2003	2003	UH357	04-AUG-2003	40.809	-73.829	1	15.2	m	
R-EMAP Region 2 2003	2003	UH357	05-AUG-2003	40.809	-73.829	2	15.2	m	
R-EMAP Region 2 2003	2003	UH358	10-JUL-2003	40.8	-73.798	1	3.0	m	
R-EMAP Region 2 2003	2003	UH358	11-JUL-2003	40.8	-73.798	2	3.0	m	
R-EMAP Region 2 2003	2003	UH359	04-AUG-2003	40.805	-73.848	1	14.9	m	
R-EMAP Region 2 2003	2003	UH359	05-AUG-2003	40.805	-73.848	2	14.9	m	
R-EMAP Region 2 2003	2003	UH360	23-AUG-2003	40.803	-73.81	1	8.5	m	
R-EMAP Region 2 2003	2003	UH360	25-AUG-2003	40.803	-73.81	2	8.5	m	
R-EMAP Region 2 2003	2003	UH361	25-AUG-2003	40.801	-73.904	1	5.8	m	
R-EMAP Region 2 2003	2003	UH361	26-AUG-2003	40.801	-73.904	2	5.8	m	
R-EMAP Region 2 2003	2003	UH361	03-SEP-2003	40.801	-73.904	3	5.8	m	
R-EMAP Region 2 2003	2003	UH362	21-JUL-2003	40.798	-73.869	1	12.5	m	
R-EMAP Region 2 2003	2003	UH363	20-AUG-2003	40.776	-73.889	1	4.0	m	
R-EMAP Region 2 2003	2003	UH363	21-AUG-2003	40.776	-73.889	2	4.0	m	
R-EMAP Region 2 2003	2003	UH365	25-AUG-2003	40.666	-74.088	1	5.2	m	
R-EMAP Region 2 2003	2003	UH365	26-AUG-2003	40.666	-74.088	2	5.2	m	
R-EMAP Region 2 2003	2003	UH366	29-AUG-2003	40.903	-73.919	1	5.2	m	
R-EMAP Region 2 2003	2003	UH366	02-SEP-2003	40.903	-73.919	2	5.2	m	
R-EMAP Region 2 2003	2003	UH366	03-SEP-2003	40.903	-73.919	3	5.2	m	
R-EMAP Region 2 2003	2003	UH368	29-AUG-2003	40.642	-74.056	1	4.9	m	
R-EMAP Region 2 2003	2003	UH368	02-SEP-2003	40.642	-74.056	2	4.9	m	
R-EMAP Region 2 2003	2003	UH369	11-SEP-2003	40.807	-73.845	1	15.2	m	
R-EMAP Region 2 2003	2003	UH369	12-SEP-2003	40.807	-73.845	2	15.2	m	
National Coastal Assessment-Southeast/Virginia Institute of Marine Sciences	2000	VA00-0001	20-SEP-2000	37.323	-77.078	1	0.9	m	
National Coastal Assessment-Southeast/Virginia Institute of Marine Sciences	2000	VA00-0002	22-SEP-2000	37.225	-76.795	1	2.1	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA00-0003	13-SEP-2001	37.325	-75.992	1	0.6	m	
National Coastal Assessment-Southeast/Virginia Institute of Marine Sciences	2000	VA00-0004	13-SEP-2000	37.696	-76.03	1	10.4	m	
National Coastal Assessment-Southeast/Virginia Institute of Marine Sciences	2000	VA00-0005	13-SEP-2000	37.611	-76.214	1	8.7	m	
National Coastal Assessment-Southeast/Virginia Institute of Marine Sciences	2000	VA00-0006	14-SEP-2000	37.542	-76.308	1	0.9	m	
National Coastal Assessment-Southeast/Virginia Institute of Marine Sciences	2000	VA00-0007	12-SEP-2000	37.331	-76.226	1	11.1	m	
National Coastal Assessment-Southeast/Virginia Institute of Marine Sciences	2000	VA00-0008	13-SEP-2000	37.722	-75.941	1	14.6	m	
National Coastal Assessment-Southeast/Virginia Institute of Marine Sciences	2000	VA00-0009	13-SEP-2000	37.615	-76.102	1	12.3	m	
National Coastal Assessment-Southeast/Virginia Institute of Marine Sciences	2000	VA00-0010	13-SEP-2000	37.567	-76.194	1	10.3	m	
National Coastal Assessment-Southeast/Virginia Institute of Marine Sciences	2000	VA00-0011	12-SEP-2000	37.463	-76.106	1	10.9	m	
National Coastal Assessment-Southeast/Virginia Institute of Marine Sciences	2000	VA00-0012	12-SEP-2000	37.224	-76.085	1	13.3	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA00-0013	27-AUG-2001	37.783	-75.803	1	0.6	m	
National Coastal Assessment-Southeast/Virginia Institute of Marine Sciences	2000	VA00-0014	13-SEP-2000	37.637	-75.925	1	5.3	m	
National Coastal Assessment-Southeast/Virginia Institute of Marine Sciences	2000	VA00-0015	12-SEP-2000	37.401	-76.041	1	12.1	m	
National Coastal Assessment-Southeast/Virginia Institute of Marine Sciences	2000	VA00-0016	12-SEP-2000	37.225	-76.035	1	6.2	m	
National Coastal Assessment-Southeast/Virginia Institute of Marine Sciences	2000	VA00-0017	11-SEP-2000	37.168	-76.011	1	8.1	m	
National Coastal Assessment-Southeast/Virginia Institute of Marine Sciences	2000	VA00-0018	11-SEP-2000	37.036	-75.975	1	5.8	m	
National Coastal Assessment-Southeast/Virginia Institute of Marine Sciences	2000	VA00-0019	12-SEP-2000	37.216	-76.27	1	5.9	m	
National Coastal Assessment-Southeast/Virginia Institute of Marine Sciences	2000	VA00-0020	11-SEP-2000	37.083	-76.16	1	10.1	m	
National Coastal Assessment-Southeast/Virginia Institute of Marine Sciences	2000	VA00-0021	11-SEP-2000	36.96	-76.008	1	19.6	m	
National Coastal Assessment-Southeast/Virginia Institute of Marine Sciences	2000	VA00-0022	27-SEP-2000	37.151	-76.244	1	8.8	m	
National Coastal Assessment-Southeast/Virginia Institute of Marine Sciences	2000	VA00-0023	27-SEP-2000	37.018	-76.258	1	4.9	m	
National Coastal Assessment-Southeast/Virginia Institute of Marine Sciences	2000	VA00-0024	20-SEP-2000	36.962	-76.401	1	2.1	m	
National Coastal Assessment-Southeast/Virginia Institute of Marine Sciences	2000	VA00-0025	27-SEP-2000	36.997	-76.254	1	5.6	m	
National Coastal Assessment-Southeast/Virginia Institute of Marine Sciences	2000	VA00-0026	11-SEP-2000	36.957	-76.098	1	9.4	m	
National Coastal Assessment-Southeast/Virginia Institute of Marine Sciences	2000	VA00-0027	15-SEP-2000	37.604	-76.367	1	8.5	m	
National Coastal Assessment-Southeast/Virginia Institute of Marine Sciences	2000	VA00-0028	18-SEP-2000	37.791	-76.649	1	1.1	m	
National Coastal Assessment-Southeast/Virginia Institute of Marine Sciences	2000	VA00-0029	18-SEP-2000	37.843	-76.751	1	2.0	m	
National Coastal Assessment-Southeast/Virginia Institute of Marine Sciences	2000	VA00-0030	18-SEP-2000	37.919	-76.831	1	0.9	m	
National Coastal Assessment-Southeast/Virginia Institute of Marine Sciences	2000	VA00-0031	07-SEP-2000	37.41	-76.674	1	1.0	m	
National Coastal Assessment-Southeast/Virginia Institute of Marine Sciences	2000	VA00-0032	07-SEP-2000	37.358	-76.634	1	2.7	m	
National Coastal Assessment-Southeast/Virginia Institute of Marine Sciences	2000	VA00-0033	08-SEP-2000	37.304	-76.579	1	3.0	m	
National Coastal Assessment-Southeast/Virginia Institute of Marine Sciences	2000	VA00-0034	20-SEP-2000	37.022	-76.503	1	2.1	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA00-0035	23-AUG-2001	36.823	-76.291	1	13.0	m	
National Coastal Assessment-Southeast/Virginia Institute of Marine Sciences	2000	VA00-0036	08-SEP-2000	37.384	-76.4	1	6.7	m	
National Coastal Assessment-Southeast/Virginia Institute of Marine Sciences	2000	VA00-0037	08-SEP-2000	37.321	-76.364	1	5.2	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0001	30-AUG-2001	37.127	-76.68	1	1.9	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0002	30-AUG-2001	37.176	-76.604	1	1.5	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0003	11-JUL-2001	37.367	-77.376	1	1.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0005	28-AUG-2001	37.3	-76.618	1	0.3	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0006	22-AUG-2001	37.331	-76.275	1	1.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0007	25-JUL-2001	37.575	-76.963	1	1.5	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0008	14-AUG-2001	37.843	-76.249	1	0.6	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0009	16-AUG-2001	37.931	-76.686	1	1.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0010	25-JUL-2001	37.79	-75.565	1	0.4	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0011	16-JUL-2001	37.616	-76.338	1	1.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0012	11-SEP-2001	38.155	-77.168	1	0.6	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0016	08-AUG-2001	36.903	-76.292	1	4.4	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0017	20-AUG-2001	36.892	-76.021	1	0.7	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0018	09-JUL-2001	36.921	-76.181	1	5.5	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0019	31-JUL-2001	37.083	-76.333	1	1.5	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0020	05-SEP-2001	37.232	-76.987	1	1.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0021	19-JUL-2001	37.109	-75.957	1	2.5	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0022	13-SEP-2001	37.44	-75.932	1	0.3	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0023	19-JUL-2001	37.616	-76.338	1	1.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0024	02-AUG-2001	37.59	-75.916	1	1.5	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0025	27-AUG-2001	37.725	-75.817	1	3.9	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0026	16-AUG-2001	37.825	-75.517	1	1.3	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0027	10-SEP-2001	37.891	-75.305	1	2.3	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0028	13-SEP-2001	38.54	-77.286	1	1.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0029	14-AUG-2001	36.836	-76.56	1	0.2	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0030	08-AUG-2001	36.848	-76.315	1	0.9	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0031	16-AUG-2001	37.309	-75.812	1	1.4	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0032	17-JUL-2001	37.562	-76.879	1	1.5	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0033	09-JUL-2001	37.538	-76.314	1	5.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0034	31-JUL-2001	37.663	-76.471	1	1.5	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0035	07-AUG-2001	37.808	-76.288	1	5.5	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0036	31-JUL-2001	37.189	-76.394	1	0.5	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0037	02-AUG-2001	37.312	-76.982	1	1.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0038	15-AUG-2001	37.579	-76.951	1	1.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0039	02-AUG-2001	37.546	-75.934	1	0.3	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0040	08-AUG-2001	37.719	-76.546	1	1.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0041	26-JUL-2001	37.922	-76.722	1	1.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0042	17-JUL-2001	36.638	-76.066	1	1.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0043	08-AUG-2001	36.84	-76.276	1	9.7	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0044	20-AUG-2001	36.871	-76.0	1	1.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0045	16-JUL-2001	37.001	-76.612	1	0.4	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0046	30-JUL-2001	37.271	-77.376	1	1.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0047	13-AUG-2001	37.358	-76.267	1	1.5	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0048	17-SEP-2001	37.338	-76.846	1	0.6	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0049	09-AUG-2001	37.568	-76.575	1	1.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2001	VA01-0050	05-JUL-2001	38.109	-76.713	1	3.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0001	09-SEP-2002	37.975	-75.405	1	1.7	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0002	17-SEP-2002	37.592	-75.633	1	2.7	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0003	03-SEP-2002	37.949	-75.422	1	0.9	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0004	16-SEP-2002	37.895	-75.454	1	2.1	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0005	19-AUG-2002	37.306	-75.806	1	0.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0006	03-SEP-2002	37.956	-75.434	1	1.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0007	15-JUL-2002	36.596	-75.913	1	0.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0008	09-SEP-2002	37.987	-75.378	1	2.1	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0009	23-SEP-2002	38.02	-75.316	1	2.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0010	15-JUL-2002	36.623	-75.942	1	0.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0011	26-AUG-2002	37.46	-75.675	1	0.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0012	23-SEP-2002	38.018	-75.281	1	0.6	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0013	26-AUG-2002	37.5	-75.734	1	0.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0014	09-SEP-2002	37.989	-75.397	1	1.9	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0015	15-JUL-2002	36.564	-75.915	1	0.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0016	29-JUL-2002	38.133	-76.645	1	1.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0017	20-AUG-2002	36.853	-76.302	1	0.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0018	16-JUL-2002	37.393	-76.25	1	0.8	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0019	01-AUG-2002	38.638	-77.208	1	1.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0020	05-AUG-2002	38.437	-77.37	1	0.8	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0021	25-JUL-2002	37.325	-76.453	1	3.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0022	18-JUL-2002	37.264	-76.877	1	7.5	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0023	17-JUL-2002	36.884	-76.016	1	1.5	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0024	29-JUL-2002	38.102	-76.732	1	1.5	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0025	30-JUL-2002	37.079	-76.305	1	0.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0026	31-JUL-2002	37.793	-75.762	1	0.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0027	15-JUL-2002	37.336	-76.28	1	1.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0029	15-AUG-2002	38.585	-77.267	1	0.6	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0030	01-AUG-2002	37.08	-76.538	1	0.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0031	30-JUL-2002	37.104	-76.32	1	4.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0032	12-AUG-2002	37.529	-76.4	1	4.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0033	07-AUG-2002	37.392	-76.413	1	0.6	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0034	08-JUL-2002	37.835	-76.281	1	4.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0035	01-AUG-2002	38.611	-77.219	1	2.5	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0036	24-JUL-2002	37.987	-76.807	1	3.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0037	18-JUL-2002	37.259	-76.872	1	5.5	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0038	08-JUL-2002	37.5	-75.91	1	0.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0039	05-AUG-2002	38.344	-77.296	1	1.5	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0040	17-JUL-2002	36.891	-76.08	1	0.7	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0041	20-AUG-2002	36.759	-76.303	1	0.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0042	19-AUG-2002	37.575	-76.978	1	1.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0043	09-JUL-2002	37.24	-76.991	1	1.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0044	01-AUG-2002	37.106	-76.682	1	0.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0045	01-JUL-2002	37.4	-76.48	1	1.2	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0046	16-JUL-2002	37.42	-76.256	1	0.4	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0047	15-AUG-2002	38.683	-77.17	1	1.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0048	02-JUL-2002	37.321	-77.28	1	2.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0049	20-AUG-2002	36.891	-76.327	1	0.0	m	
National Coastal Assessment-Southeast/Virginia Department of Environmental Quality	2002	VA02-0050	07-AUG-2002	37.43	-76.452	1	3.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0001-A	25-JUL-2005	37.378	-76.898	1	0.6	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0001-A	31-AUG-2005	37.378	-76.898	1	0.6	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0002-A	01-AUG-2005	37.191	-76.106	1	9.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0002-A	09-SEP-2005	37.191	-76.106	2	9.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0003-A	30-AUG-2005	37.059	-76.595	1	4.2	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0003-A	20-SEP-2005	37.059	-76.595	2	4.2	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0004-A	25-JUL-2005	37.579	-76.964	1	0.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0004-A	31-AUG-2005	37.579	-76.964	1	0.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0006-A	06-JUL-2005	37.649	-76.486	1	7.4	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0007-A	12-JUL-2005	37.322	-77.196	1	1.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0008-A	01-SEP-2005	37.28	-76.544	1	5.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0008-A	08-SEP-2005	37.28	-76.544	2	5.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0009-A	09-AUG-2005	36.911	-76.461	1	2.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0010-A	01-AUG-2005	37.248	-76.13	1	14.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0010-A	09-SEP-2005	37.248	-76.13	2	14.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0011-A	02-AUG-2005	37.59	-76.195	1	12.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0011-A	13-SEP-2005	37.59	-76.195	2	12.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0012-A	14-JUL-2005	37.979	-75.345	1	1.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0013-A	20-JUL-2005	37.673	-75.855	1	2.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0014-A	19-JUL-2005	37.763	-75.769	1	3.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0015-A	02-AUG-2005	37.446	-76.087	1	16.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0015-A	12-SEP-2005	37.446	-76.087	2	16.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0016-A	14-JUL-2005	37.947	-76.867	1	1.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0017-A	07-JUL-2005	36.83	-76.393	1	2.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0018-B	01-AUG-2005	37.091	-76.009	1	6.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0018-B	19-SEP-2005	37.091	-76.009	2	6.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0019-A	28-JUL-2005	36.996	-76.495	1	4.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0020-A	19-JUL-2005	37.466	-76.746	1	1.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0021-A	01-AUG-2005	37.003	-76.005	1	9.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0021-A	19-SEP-2005	37.003	-76.005	2	9.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0022-A	26-JUL-2005	37.612	-76.509	1	1.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0022-A	16-SEP-2005	37.612	-76.509	2	1.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0023-A	21-JUL-2005	37.283	-77.081	1	9.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0024-A	01-AUG-2005	37.013	-76.285	1	7.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0024-A	22-SEP-2005	37.013	-76.285	2	7.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0025-A	02-AUG-2005	37.714	-76.035	1	10.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0025-A	13-SEP-2005	37.714	-76.035	2	10.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0026-A	22-JUL-2005	37.375	-76.454	1	1.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0026-A	08-SEP-2005	37.375	-76.454	1	1.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0027-A	15-AUG-2005	37.628	-76.398	1	6.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0028-A	14-JUL-2005	38.012	-75.368	1	2.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0028-A	22-AUG-2005	38.012	-75.368	2	2.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0029-A	26-JUL-2005	37.703	-76.461	1	4.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0029-A	16-SEP-2005	37.703	-76.461	1	4.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0030-A	24-AUG-2005	37.891	-75.793	1	4.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0030-A	07-SEP-2005	37.891	-75.793	1	4.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0031-A	04-AUG-2005	37.313	-75.822	1	0.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0031-A	24-AUG-2005	37.313	-75.822	2	0.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0032-A	26-JUL-2005	38.145	-77.05	1	1.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0033-A	12-JUL-2005	36.948	-76.404	1	8.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0034-A	26-JUL-2005	37.169	-75.921	1	1.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0035-A	17-AUG-2005	37.795	-76.315	1	1.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0036-B	11-AUG-2005	37.904	-75.469	1	1.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0036-B	22-AUG-2005	37.904	-75.469	2	1.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0037-A	02-AUG-2005	37.776	-76.073	1	7.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0037-A	13-SEP-2005	37.776	-76.073	2	7.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0038-A	02-AUG-2005	37.89	-75.409	1	2.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0038-A	22-AUG-2005	37.89	-75.409	2	2.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0039-A	04-AUG-2005	37.333	-75.796	1	1.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0039-A	24-AUG-2005	37.333	-75.796	2	1.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0040-A	11-AUG-2005	37.841	-76.759	1	1.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0041-A	27-JUL-2005	36.876	-76.059	1	0.6	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0041-A	30-AUG-2005	36.876	-76.059	1	0.6	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0042-A	11-AUG-2005	37.776	-76.666	1	6.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0043-A	02-AUG-2005	37.13	-76.652	1	5.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0044-A	27-JUL-2005	37.254	-76.43	1	0.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0044-A	01-SEP-2005	37.254	-76.43	1	0.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0046-A	22-JUL-2005	37.526	-76.436	1	1.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0046-A	08-SEP-2005	37.526	-76.436	1	1.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0047-A	04-AUG-2005	37.189	-76.773	1	5.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0048-A	25-AUG-2005	37.16	-76.393	1	1.4	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0049-A	12-JUL-2005	36.927	-76.411	1	5.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0050-A	16-SEP-2005	37.785	-76.641	1	2.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2005	VA05-0050-A	18-SEP-2005	37.785	-76.641	1	2.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0051-A	17-AUG-2006	36.953	-76.277	1	3.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0052-B	03-AUG-2006	37.195	-75.864	1	1.7	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0052-B	29-AUG-2006	37.195	-75.864	1	5.2	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0053-A	19-JUL-2006	37.754	-76.254	1	7.1	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0053-A	25-SEP-2006	37.754	-76.254	1	6.7	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0054-A	26-JUL-2006	37.95	-75.407	1	4.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0055-A	07-SEP-2006	37.729	-75.845	1	1.4	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0055-A	18-SEP-2006	37.729	-75.845	1	1.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0056-A	27-JUL-2006	37.623	-75.657	1	0.7	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0056-A	24-AUG-2006	37.623	-75.657	1	4.3	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0057-C	28-SEP-2006	37.48	-75.807	1	3.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0058-A	19-JUL-2006	37.881	-76.146	1	20.3	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0058-A	25-SEP-2006	37.881	-76.146	1	20.4	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0059-A	18-JUL-2006	36.875	-76.332	1	15.6	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0059-A	31-JUL-2006	36.875	-76.332	1	2.4	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0060-A	25-JUL-2006	37.75	-76.635	1	1.2	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0060-A	06-SEP-2006	37.75	-76.635	1	0.9	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0061-A	21-SEP-2006	37.063	-76.67	1	1.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0062-A	13-JUL-2006	37.353	-76.633	1	4.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0064-A	10-AUG-2006	37.617	-76.477	1	5.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0065-A	18-JUL-2006	37.218	-76.895	1	3.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0066-A	08-AUG-2006	37.024	-76.497	1	2.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0067-A	18-JUL-2006	36.999	-76.342	1	3.8	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0067-A	31-JUL-2006	36.999	-76.342	1	4.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0068-A	03-AUG-2006	37.137	-75.938	1	1.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0069-A	19-JUL-2006	37.518	-76.055	1	14.8	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0069-A	22-SEP-2006	37.518	-76.055	1	14.6	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0070-A	02-AUG-2006	37.929	-75.343	1	1.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0071-A	19-JUL-2006	37.576	-75.989	1	11.8	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0071-A	22-SEP-2006	37.576	-75.989	1	11.3	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0072-B	24-AUG-2006	37.891	-75.405	1	0.9	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0072-B	20-SEP-2006	37.891	-75.405	1	5.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0073-A	20-JUL-2006	37.328	-76.021	1	3.3	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0073-A	18-SEP-2006	37.328	-76.021	1	3.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0074-A	19-JUL-2006	37.914	-76.8	1	1.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0076-A	06-SEP-2006	37.635	-76.522	1	14.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0076-A	25-SEP-2006	37.635	-76.522	1	13.7	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0077-A	31-JUL-2006	37.182	-76.696	1	1.2	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0077-A	09-AUG-2006	37.182	-76.696	1	1.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0078-A	25-JUL-2006	37.23	-76.492	1	7.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0080-A	24-JUL-2006	37.487	-76.347	1	1.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0080-A	13-SEP-2006	37.487	-76.347	1	0.9	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0081-A	26-JUL-2006	37.266	-76.881	1	3.4	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0081-A	09-AUG-2006	37.266	-76.881	1	3.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0082-A	05-SEP-2006	37.113	-76.566	1	4.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0083-A	27-JUL-2006	37.358	-77.304	1	4.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0084-A	18-JUL-2006	37.069	-76.122	1	10.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0084-A	08-SEP-2006	37.069	-76.122	1	11.9	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0085-A	25-JUL-2006	37.005	-76.582	1	1.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0086-A	01-AUG-2006	37.402	-76.676	1	6.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0088-A	08-AUG-2006	37.703	-76.554	1	10.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0089-A	26-JUL-2006	37.311	-77.304	1	4.3	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0089-A	10-AUG-2006	37.311	-77.304	1	5.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0090-A	02-AUG-2006	37.094	-76.347	1	2.7	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0090-A	11-SEP-2006	37.094	-76.347	1	1.1	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0091-A	11-JUL-2006	36.762	-76.307	1	2.5	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0092-A	18-JUL-2006	37.34	-76.335	1	4.4	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0092-A	24-JUL-2006	37.34	-76.335	1	3.7	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0093-A	15-AUG-2006	37.522	-76.31	1	6.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0094-A	26-JUL-2006	38.012	-75.312	1	1.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0095-A	20-JUL-2006	37.505	-75.7	1	2.4	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0096-C	07-SEP-2006	37.699	-75.611	1	4.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0097-A	13-JUL-2006	37.33	-75.891	1	4.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0097-A	29-AUG-2006	37.33	-75.891	1	4.3	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0098-A	25-JUL-2006	38.108	-77.003	1	0.9	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0098-A	12-SEP-2006	38.108	-77.003	1	0.9	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0099-A	25-SEP-2006	36.982	-76.478	1	3.0	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0100-A	18-JUL-2006	37.254	-76.249	1	10.2	m	
National Coastal Assessment-Northeast/USEPA Office of Research and Development	2006	VA06-0100-A	13-SEP-2006	37.254	-76.249	1	9.4	m	
EMAP Virginian Province	1990	VA90-001	29-AUG-1990	38.862	-75.109	1	22.7	m	
EMAP Virginian Province	1990	VA90-002	29-AUG-1990	39.155	-74.925	1			
EMAP Virginian Province	1990	VA90-003	29-AUG-1990	39.149	-75.031	1			
EMAP Virginian Province	1990	VA90-004	29-AUG-1990	39.145	-75.135	1	3.5	m	
EMAP Virginian Province	1990	VA90-005	24-JUL-1990	39.138	-75.254	1	9.1	m	
EMAP Virginian Province	1990	VA90-006	24-JUL-1990	39.133	-75.34	1	4.9	m	
EMAP Virginian Province	1990	VA90-007	24-JUL-1990	39.204	-75.295	1	7.2	m	
EMAP Virginian Province	1990	VA90-008	31-AUG-1990	39.277	-75.25	1	3.9	m	
EMAP Virginian Province	1990	VA90-009	31-AUG-1990	39.27	-75.372	1			
EMAP Virginian Province	1990	VA90-010	30-AUG-1990	39.337	-75.438	1	8.7	m	
EMAP Virginian Province	1990	VA90-011	30-AUG-1990	39.464	-75.562	1			
EMAP Virginian Province	1990	VA90-012	04-AUG-1990	38.856	-75.216	1	3.6	m	
EMAP Virginian Province	1990	VA90-012	28-AUG-1990	38.856	-75.216	2			
EMAP Virginian Province	1990	VA90-013	30-AUG-1990	39.404	-75.491	1	7.8	m	
EMAP Virginian Province	1990	VA90-014	28-AUG-1990	38.939	-75.067	1	9.9	m	
EMAP Virginian Province	1990	VA90-015	28-AUG-1990	38.925	-75.28	1	3.4	m	
EMAP Virginian Province	1990	VA90-016	29-AUG-1990	39.012	-75.025	1			
EMAP Virginian Province	1990	VA90-017	28-AUG-1990	39.005	-75.133	1	6.7	m	
EMAP Virginian Province	1990	VA90-018	03-AUG-1990	38.999	-75.232	1	16.9	m	
EMAP Virginian Province	1990	VA90-019	29-AUG-1990	39.083	-74.986	1	5.6	m	
EMAP Virginian Province	1990	VA90-020	03-AUG-1990	39.069	-75.196	1	8.5	m	
EMAP Virginian Province	1990	VA90-021	21-JUL-1990	41.03	-72.804	1	39.0	m	
EMAP Virginian Province	1990	VA90-021	13-SEP-1990	41.03	-72.804	2	38.8	m	
EMAP Virginian Province	1990	VA90-022	23-JUL-1990	41.166	-72.926	1	16.5	m	
EMAP Virginian Province	1990	VA90-022	01-AUG-1990	41.166	-72.926	2	17.0	m	
EMAP Virginian Province	1990	VA90-022	13-AUG-1990	41.166	-72.926	3	16.6	m	
EMAP Virginian Province	1990	VA90-022	22-AUG-1990	41.166	-72.926	4	16.8	m	
EMAP Virginian Province	1990	VA90-022	30-AUG-1990	41.166	-72.926	5	16.7	m	
EMAP Virginian Province	1990	VA90-022	14-SEP-1990	41.166	-72.926	6	18.2	m	
EMAP Virginian Province	1990	VA90-023	19-AUG-1990	40.741	-72.998	1	2.2	m	
EMAP Virginian Province	1990	VA90-023	28-AUG-1990	40.741	-72.998	2	2.0	m	
EMAP Virginian Province	1990	VA90-023	12-SEP-1990	40.741	-72.998	3	2.2	m	
EMAP Virginian Province	1990	VA90-024	21-JUL-1990	41.021	-73.023	1	40.9	m	
EMAP Virginian Province	1990	VA90-024	13-SEP-1990	41.021	-73.023	2	41.3	m	
EMAP Virginian Province	1990	VA90-025	22-JUL-1990	41.012	-73.242	1	36.7	m	
EMAP Virginian Province	1990	VA90-025	23-SEP-1990	41.012	-73.242	2	34.0	m	
EMAP Virginian Province	1990	VA90-026	22-JUL-1990	41.002	-73.461	1	24.0	m	
EMAP Virginian Province	1990	VA90-026	01-AUG-1990	41.002	-73.461	2	27.5	m	
EMAP Virginian Province	1990	VA90-026	09-AUG-1990	41.002	-73.461	3	25.3	m	
EMAP Virginian Province	1990	VA90-026	29-AUG-1990	41.002	-73.461	4	26.4	m	
EMAP Virginian Province	1990	VA90-026	22-SEP-1990	41.002	-73.461	5	27.6	m	
EMAP Virginian Province	1990	VA90-027	05-AUG-1990	41.525	-70.072	1	5.6	m	
EMAP Virginian Province	1990	VA90-027	27-SEP-1990	41.525	-70.072	2	5.6	m	
EMAP Virginian Province	1990	VA90-028	31-JUL-1990	40.846	-73.775	1	6.2	m	
EMAP Virginian Province	1990	VA90-028	22-SEP-1990	40.846	-73.775	2	7.1	m	
EMAP Virginian Province	1990	VA90-029	05-AUG-1990	41.383	-70.177	1	12.8	m	
EMAP Virginian Province	1990	VA90-029	27-SEP-1990	41.383	-70.177	2	12.5	m	
EMAP Virginian Province	1990	VA90-031	29-AUG-1990	39.077	-75.088	1			
EMAP Virginian Province	1990	VA90-031	12-SEP-1990	39.077	-75.088	2	7.3	m	
EMAP Virginian Province	1990	VA90-032	04-AUG-1990	38.929	-75.176	1	15.3	m	
EMAP Virginian Province	1990	VA90-032	12-SEP-1990	38.929	-75.176	2			
EMAP Virginian Province	1990	VA90-033	23-JUL-1990	39.21	-75.212	1	4.4	m	
EMAP Virginian Province	1990	VA90-033	03-AUG-1990	39.21	-75.212	2	6.2	m	
EMAP Virginian Province	1990	VA90-033	12-AUG-1990	39.21	-75.212	3	5.0	m	
EMAP Virginian Province	1990	VA90-033	22-AUG-1990	39.21	-75.212	4	7.2	m	
EMAP Virginian Province	1990	VA90-033	30-AUG-1990	39.21	-75.212	5	6.6	m	
EMAP Virginian Province	1990	VA90-033	12-SEP-1990	39.21	-75.212	6	5.6	m	
EMAP Virginian Province	1990	VA90-034	18-AUG-1990	38.073	-75.275	1	2.0	m	
EMAP Virginian Province	1990	VA90-034	17-SEP-1990	38.073	-75.275	2	2.4	m	
EMAP Virginian Province	1990	VA90-035	03-AUG-1990	39.063	-75.3	1	5.1	m	
EMAP Virginian Province	1990	VA90-035	12-SEP-1990	39.063	-75.3	2	4.6	m	
EMAP Virginian Province	1990	VA90-036	31-AUG-1990	39.343	-75.337	1	2.4	m	
EMAP Virginian Province	1990	VA90-036	09-SEP-1990	39.343	-75.337	2	3.4	m	
EMAP Virginian Province	1990	VA90-037	16-AUG-1990	41.522	-70.294	1	10.6	m	
EMAP Virginian Province	1990	VA90-037	06-SEP-1990	41.522	-70.294	2	11.2	m	
EMAP Virginian Province	1990	VA90-038	16-AUG-1990	41.38	-70.398	1	14.4	m	
EMAP Virginian Province	1990	VA90-038	06-SEP-1990	41.38	-70.398	2	13.0	m	
EMAP Virginian Province	1990	VA90-039	11-AUG-1990	37.895	-75.778	1	4.0	m	
EMAP Virginian Province	1990	VA90-040	19-AUG-1990	37.747	-75.862	1	7.0	m	
EMAP Virginian Province	1990	VA90-040	16-SEP-1990	37.747	-75.862	2	5.5	m	
EMAP Virginian Province	1990	VA90-041	20-JUL-1990	38.028	-75.902	1	4.9	m	
EMAP Virginian Province	1990	VA90-041	29-JUL-1990	38.028	-75.902	2	5.1	m	
EMAP Virginian Province	1990	VA90-041	08-AUG-1990	38.028	-75.902	3	5.4	m	
EMAP Virginian Province	1990	VA90-041	19-AUG-1990	38.028	-75.902	4	5.3	m	
EMAP Virginian Province	1990	VA90-041	29-AUG-1990	38.028	-75.902	5	5.2	m	
EMAP Virginian Province	1990	VA90-041	18-SEP-1990	38.028	-75.902	6	6.1	m	
EMAP Virginian Province	1990	VA90-042	03-AUG-1990	37.599	-75.945	1			
EMAP Virginian Province	1990	VA90-042	05-SEP-1990	37.599	-75.945	2	7.2	m	
EMAP Virginian Province	1990	VA90-044	21-JUL-1990	37.17	-75.988	1	5.7	m	
EMAP Virginian Province	1990	VA90-045	20-JUL-1990	38.16	-76.026	1	1.5	m	
EMAP Virginian Province	1990	VA90-045	20-SEP-1990	38.16	-76.026	2			
EMAP Virginian Province	1990	VA90-046	04-AUG-1990	37.45	-76.028	1	14.2	m	
EMAP Virginian Province	1990	VA90-046	05-SEP-1990	37.45	-76.028	2			
EMAP Virginian Province	1990	VA90-047	29-JUL-1990	37.731	-76.069	1			
EMAP Virginian Province	1990	VA90-047	16-SEP-1990	37.731	-76.069	2	9.1	m	
EMAP Virginian Province	1990	VA90-048	22-JUL-1990	37.021	-76.07	1	13.8	m	
EMAP Virginian Province	1990	VA90-048	12-SEP-1990	37.021	-76.07	2	10.0	m	
EMAP Virginian Province	1990	VA90-050	20-JUL-1990	38.012	-76.11	1	7.7	m	
EMAP Virginian Province	1990	VA90-050	20-SEP-1990	38.012	-76.11	2			
EMAP Virginian Province	1990	VA90-051	31-JUL-1990	37.302	-76.111	1	17.6	m	
EMAP Virginian Province	1990	VA90-052	26-AUG-1990	41.518	-70.516	1	2.4	m	
EMAP Virginian Province	1990	VA90-052	05-SEP-1990	41.518	-70.516	2	2.5	m	
EMAP Virginian Province	1990	VA90-053	03-AUG-1990	37.583	-76.153	1			
EMAP Virginian Province	1990	VA90-053	05-SEP-1990	37.583	-76.153	2			
EMAP Virginian Province	1990	VA90-054	21-JUL-1990	37.153	-76.193	1	10.6	m	
EMAP Virginian Province	1990	VA90-054	31-JUL-1990	37.153	-76.193	2	10.7	m	
EMAP Virginian Province	1990	VA90-054	09-AUG-1990	37.153	-76.193	3	10.9	m	
EMAP Virginian Province	1990	VA90-054	20-AUG-1990	37.153	-76.193	4	10.5	m	
EMAP Virginian Province	1990	VA90-054	29-AUG-1990	37.153	-76.193	5	11.3	m	
EMAP Virginian Province	1990	VA90-055	24-AUG-1990	37.864	-76.194	1	8.9	m	
EMAP Virginian Province	1990	VA90-055	16-SEP-1990	37.864	-76.194	2	9.5	m	
EMAP Virginian Province	1990	VA90-056	19-AUG-1990	38.144	-76.235	1	14.4	m	
EMAP Virginian Province	1990	VA90-057	25-JUL-1990	37.434	-76.235	1	2.4	m	
EMAP Virginian Province	1990	VA90-057	06-SEP-1990	37.434	-76.235	2	2.5	m	
EMAP Virginian Province	1990	VA90-058	17-AUG-1990	39.129	-76.281	1	2.2	m	
EMAP Virginian Province	1990	VA90-058	08-SEP-1990	39.129	-76.281	2			
EMAP Virginian Province	1990	VA90-059	22-JUL-1990	37.005	-76.275	1	11.2	m	
EMAP Virginian Province	1990	VA90-059	12-SEP-1990	37.005	-76.275	2	10.0	m	
EMAP Virginian Province	1990	VA90-060	03-AUG-1990	37.715	-76.277	1	6.6	m	
EMAP Virginian Province	1990	VA90-060	05-SEP-1990	37.715	-76.277	2			
EMAP Virginian Province	1990	VA90-061	25-JUL-1990	37.286	-76.318	1	7.9	m	
EMAP Virginian Province	1990	VA90-061	04-AUG-1990	37.286	-76.318	2	7.3	m	
EMAP Virginian Province	1990	VA90-061	13-AUG-1990	37.286	-76.318	3	8.2	m	
EMAP Virginian Province	1990	VA90-061	23-AUG-1990	37.286	-76.318	4	8.5	m	
EMAP Virginian Province	1990	VA90-061	06-SEP-1990	37.286	-76.318	5	8.6	m	
EMAP Virginian Province	1990	VA90-062	24-AUG-1990	38.987	-76.358	1	25.5	m	
EMAP Virginian Province	1990	VA90-062	07-SEP-1990	38.987	-76.358	2	15.7	m	
EMAP Virginian Province	1990	VA90-063	25-AUG-1990	38.277	-76.36	1	9.9	m	
EMAP Virginian Province	1990	VA90-065	27-JUL-1990	38.558	-76.401	1	8.6	m	
EMAP Virginian Province	1990	VA90-065	06-AUG-1990	38.558	-76.401	2	8.4	m	
EMAP Virginian Province	1990	VA90-065	16-AUG-1990	38.558	-76.401	3	8.8	m	
EMAP Virginian Province	1990	VA90-065	28-AUG-1990	38.558	-76.401	4	7.5	m	
EMAP Virginian Province	1990	VA90-065	07-SEP-1990	38.558	-76.401	5	8.3	m	
EMAP Virginian Province	1990	VA90-066	24-AUG-1990	38.838	-76.443	1			
EMAP Virginian Province	1990	VA90-066	04-SEP-1990	38.838	-76.443	2			
EMAP Virginian Province	1990	VA90-068	06-AUG-1990	41.371	-70.841	1	27.1	m	
EMAP Virginian Province	1990	VA90-069	26-JUL-1990	41.509	-70.959	1	7.0	m	
EMAP Virginian Province	1990	VA90-069	25-SEP-1990	41.509	-70.959	2	7.6	m	
EMAP Virginian Province	1990	VA90-070	28-JUL-1990	41.641	-71.3	1	8.9	m	
EMAP Virginian Province	1990	VA90-070	07-AUG-1990	41.641	-71.3	2	10.0	m	
EMAP Virginian Province	1990	VA90-070	17-AUG-1990	41.641	-71.3	3	10.2	m	
EMAP Virginian Province	1990	VA90-070	27-AUG-1990	41.641	-71.3	4	9.7	m	
EMAP Virginian Province	1990	VA90-070	08-SEP-1990	41.641	-71.3	5	9.8	m	
EMAP Virginian Province	1990	VA90-071	24-SEP-1990	41.498	-71.402	1	9.2	m	
EMAP Virginian Province	1990	VA90-072	04-AUG-1990	41.355	-71.504	1	8.4	m	
EMAP Virginian Province	1990	VA90-072	17-SEP-1990	41.355	-71.504	2	8.3	m	
EMAP Virginian Province	1990	VA90-073	04-AUG-1990	41.212	-71.605	1	32.0	m	
EMAP Virginian Province	1990	VA90-073	16-SEP-1990	41.212	-71.605	2	31.0	m	
EMAP Virginian Province	1990	VA90-074	03-AUG-1990	41.205	-71.825	1	35.1	m	
EMAP Virginian Province	1990	VA90-074	16-SEP-1990	41.205	-71.825	2	35.4	m	
EMAP Virginian Province	1990	VA90-075	03-AUG-1990	41.198	-72.046	1	48.6	m	
EMAP Virginian Province	1990	VA90-075	16-SEP-1990	41.198	-72.046	2	49.6	m	
EMAP Virginian Province	1990	VA90-076	29-JUL-1990	41.191	-72.266	1	42.7	m	
EMAP Virginian Province	1990	VA90-076	11-SEP-1990	41.191	-72.266	2	42.6	m	
EMAP Virginian Province	1990	VA90-077	13-AUG-1990	41.183	-72.486	1	12.2	m	
EMAP Virginian Province	1990	VA90-077	27-SEP-1990	41.183	-72.486	2	8.0	m	
EMAP Virginian Province	1990	VA90-078	18-AUG-1990	41.039	-72.584	1	17.8	m	
EMAP Virginian Province	1990	VA90-078	12-SEP-1990	41.039	-72.584	2	19.0	m	
EMAP Virginian Province	1990	VA90-079	13-AUG-1990	41.175	-72.706	1	26.2	m	
EMAP Virginian Province	1990	VA90-080	16-AUG-1990	38.89	-76.401	1			
EMAP Virginian Province	1990	VA90-080	07-SEP-1990	38.89	-76.401	2	21.1	m	
EMAP Virginian Province	1990	VA90-081	27-AUG-1990	39.243	-76.492	1			
EMAP Virginian Province	1990	VA90-081	06-SEP-1990	39.243	-76.492	2			
EMAP Virginian Province	1990	VA90-082	27-AUG-1990	39.253	-76.552	1			
EMAP Virginian Province	1990	VA90-082	06-SEP-1990	39.253	-76.552	2	5.5	m	
EMAP Virginian Province	1990	VA90-083	24-AUG-1990	38.878	-76.515	1	3.8	m	
EMAP Virginian Province	1990	VA90-083	04-SEP-1990	38.878	-76.515	2			
EMAP Virginian Province	1990	VA90-084	14-AUG-1990	37.623	-76.465	1	6.6	m	
EMAP Virginian Province	1990	VA90-084	07-SEP-1990	37.623	-76.465	2			
EMAP Virginian Province	1990	VA90-085	13-AUG-1990	37.067	-76.167	1			
EMAP Virginian Province	1990	VA90-085	12-SEP-1990	37.067	-76.167	2	7.5	m	
EMAP Virginian Province	1990	VA90-086	22-JUL-1990	36.832	-76.294	1	6.6	m	
EMAP Virginian Province	1990	VA90-086	01-AUG-1990	36.832	-76.294	2	5.9	m	
EMAP Virginian Province	1990	VA90-086	12-AUG-1990	36.832	-76.294	3	6.3	m	
EMAP Virginian Province	1990	VA90-086	20-AUG-1990	36.832	-76.294	4	7.0	m	
EMAP Virginian Province	1990	VA90-086	30-AUG-1990	36.832	-76.294	5	7.0	m	
EMAP Virginian Province	1990	VA90-086	13-SEP-1990	36.832	-76.294	6	7.2	m	
EMAP Virginian Province	1990	VA90-087	20-AUG-1990	37.0	-76.333	1	3.3	m	
EMAP Virginian Province	1990	VA90-087	11-SEP-1990	37.0	-76.333	2	2.5	m	
EMAP Virginian Province	1990	VA90-088	28-JUL-1990	38.87	-76.998	1	4.8	m	
EMAP Virginian Province	1990	VA90-088	07-AUG-1990	38.87	-76.998	2	6.8	m	
EMAP Virginian Province	1990	VA90-088	17-AUG-1990	38.87	-76.998	3	4.6	m	
EMAP Virginian Province	1990	VA90-088	26-AUG-1990	38.87	-76.998	4	4.9	m	
EMAP Virginian Province	1990	VA90-088	21-SEP-1990	38.87	-76.998	5			
EMAP Virginian Province	1990	VA90-089	07-AUG-1990	39.378	-76.0	1			
EMAP Virginian Province	1990	VA90-089	16-SEP-1990	39.378	-76.0	2			
EMAP Virginian Province	1990	VA90-090	26-JUL-1990	39.27	-76.443	1	1.7	m	
EMAP Virginian Province	1990	VA90-090	04-AUG-1990	39.27	-76.443	2	1.8	m	
EMAP Virginian Province	1990	VA90-090	15-AUG-1990	39.27	-76.443	3	1.7	m	
EMAP Virginian Province	1990	VA90-090	23-AUG-1990	39.27	-76.443	4	2.0	m	
EMAP Virginian Province	1990	VA90-090	05-SEP-1990	39.27	-76.443	5	2.5	m	
EMAP Virginian Province	1990	VA90-091	14-AUG-1990	39.443	-76.246	1	2.0	m	
EMAP Virginian Province	1990	VA90-091	14-SEP-1990	39.443	-76.246	2			
EMAP Virginian Province	1990	VA90-093	23-AUG-1990	41.347	-72.378	1	7.0	m	
EMAP Virginian Province	1990	VA90-093	17-SEP-1990	41.347	-72.378	2	6.1	m	
EMAP Virginian Province	1990	VA90-094	30-JUL-1990	40.622	-74.203	1	12.9	m	
EMAP Virginian Province	1990	VA90-094	20-SEP-1990	40.622	-74.203	2	4.7	m	
EMAP Virginian Province	1990	VA90-095	02-AUG-1990	41.313	-72.886	1	5.6	m	
EMAP Virginian Province	1990	VA90-095	30-AUG-1990	41.313	-72.886	2	5.6	m	
EMAP Virginian Province	1990	VA90-096	31-JUL-1990	40.92	-73.645	1	18.5	m	
EMAP Virginian Province	1990	VA90-096	21-SEP-1990	40.92	-73.645	2	19.1	m	
EMAP Virginian Province	1990	VA90-098	20-AUG-1990	41.16	-73.21	1	8.3	m	
EMAP Virginian Province	1990	VA90-098	23-SEP-1990	41.16	-73.21	2	6.9	m	
EMAP Virginian Province	1990	VA90-099	26-JUL-1990	41.643	-70.912	1	10.0	m	
EMAP Virginian Province	1990	VA90-099	06-AUG-1990	41.643	-70.912	2	10.2	m	
EMAP Virginian Province	1990	VA90-099	15-AUG-1990	41.643	-70.912	3	10.3	m	
EMAP Virginian Province	1990	VA90-099	25-AUG-1990	41.643	-70.912	5	10.7	m	
EMAP Virginian Province	1990	VA90-099	04-SEP-1990	41.643	-70.912	6	2.6	m	
EMAP Virginian Province	1990	VA90-100	21-JUL-1990	40.343	-73.987	1	2.1	m	
EMAP Virginian Province	1990	VA90-100	01-AUG-1990	40.343	-73.987	2	2.1	m	
EMAP Virginian Province	1990	VA90-100	09-AUG-1990	40.343	-73.987	3			
EMAP Virginian Province	1990	VA90-100	21-AUG-1990	40.343	-73.987	4	1.6	m	
EMAP Virginian Province	1990	VA90-100	27-AUG-1990	40.343	-73.987	5	2.0	m	
EMAP Virginian Province	1990	VA90-100	21-SEP-1990	40.343	-73.987	6			
EMAP Virginian Province	1990	VA90-101	11-AUG-1990	41.383	-73.956	1	15.0	m	
EMAP Virginian Province	1990	VA90-101	20-SEP-1990	41.383	-73.956	2	18.0	m	
EMAP Virginian Province	1990	VA90-102	01-AUG-1990	40.75	-74.087	1	5.7	m	
EMAP Virginian Province	1990	VA90-102	19-SEP-1990	40.75	-74.087	2	2.9	m	
EMAP Virginian Province	1990	VA90-103	31-JUL-1990	40.75	-74.165	1	5.8	m	
EMAP Virginian Province	1990	VA90-103	20-SEP-1990	40.75	-74.165	2	5.2	m	
EMAP Virginian Province	1990	VA90-104	20-JUL-1990	40.957	-72.503	1	6.3	m	
EMAP Virginian Province	1990	VA90-104	30-JUL-1990	40.957	-72.503	2	6.4	m	
EMAP Virginian Province	1990	VA90-104	08-AUG-1990	40.957	-72.503	3	6.2	m	
EMAP Virginian Province	1990	VA90-104	19-AUG-1990	40.957	-72.503	4	6.2	m	
EMAP Virginian Province	1990	VA90-104	28-AUG-1990	40.957	-72.503	5	6.7	m	
EMAP Virginian Province	1990	VA90-104	09-SEP-1990	40.957	-72.503	6	6.4	m	
EMAP Virginian Province	1990	VA90-105	08-AUG-1990	40.931	-72.518	1	6.3	m	
EMAP Virginian Province	1990	VA90-106	25-JUL-1990	41.365	-71.964	1	3.0	m	
EMAP Virginian Province	1990	VA90-106	03-AUG-1990	41.365	-71.964	2	2.5	m	
EMAP Virginian Province	1990	VA90-106	14-AUG-1990	41.365	-71.964	3	2.9	m	
EMAP Virginian Province	1990	VA90-106	24-AUG-1990	41.365	-71.964	4	2.6	m	
EMAP Virginian Province	1990	VA90-106	15-SEP-1990	41.365	-71.964	5	2.6	m	
EMAP Virginian Province	1990	VA90-107	14-AUG-1990	41.325	-71.977	1	2.3	m	
EMAP Virginian Province	1990	VA90-108	24-AUG-1990	41.338	-71.975	1	4.5	m	
EMAP Virginian Province	1990	VA90-111	09-AUG-1990	40.343	-74.0	1			
EMAP Virginian Province	1990	VA90-112	27-JUL-1990	38.878	-76.518	1	3.4	m	
EMAP Virginian Province	1990	VA90-112	04-SEP-1990	38.878	-76.518	2			
EMAP Virginian Province	1990	VA90-113	27-JUL-1990	38.854	-76.518	1	3.9	m	
EMAP Virginian Province	1990	VA90-114	06-AUG-1990	38.745	-76.242	1	3.6	m	
EMAP Virginian Province	1990	VA90-114	07-SEP-1990	38.745	-76.242	2	6.5	m	
EMAP Virginian Province	1990	VA90-115	06-AUG-1990	38.743	-76.242	1	6.1	m	
EMAP Virginian Province	1990	VA90-118	11-AUG-1990	39.542	-74.408	1	4.2	m	
EMAP Virginian Province	1990	VA90-118	23-SEP-1990	39.542	-74.408	2	6.1	m	
EMAP Virginian Province	1990	VA90-119	11-AUG-1990	39.518	-74.412	1	2.6	m	
EMAP Virginian Province	1990	VA90-120	11-AUG-1990	39.552	-74.415	1	2.3	m	
EMAP Virginian Province	1990	VA90-122	21-JUL-1990	40.46	-74.075	1	6.1	m	
EMAP Virginian Province	1990	VA90-122	21-SEP-1990	40.46	-74.075	2	6.5	m	
EMAP Virginian Province	1990	VA90-123	21-JUL-1990	40.442	-74.027	1			
EMAP Virginian Province	1990	VA90-124	27-AUG-1990	39.502	-75.533	1	3.1	m	
EMAP Virginian Province	1990	VA90-124	16-SEP-1990	39.502	-75.533	2	3.3	m	
EMAP Virginian Province	1990	VA90-125	27-AUG-1990	39.503	-75.534	1	3.1	m	
EMAP Virginian Province	1990	VA90-128	27-JUL-1990	38.458	-77.039	1	2.6	m	
EMAP Virginian Province	1990	VA90-128	14-SEP-1990	38.458	-77.039	2			
EMAP Virginian Province	1990	VA90-129	27-JUL-1990	38.417	-77.026	1			
EMAP Virginian Province	1990	VA90-130	11-AUG-1990	37.998	-75.622	1	4.6	m	
EMAP Virginian Province	1990	VA90-130	24-SEP-1990	37.998	-75.622	2	4.8	m	
EMAP Virginian Province	1990	VA90-132	26-JUL-1990	41.642	-70.921	1	9.3	m	
EMAP Virginian Province	1990	VA90-133	11-AUG-1990	37.963	-75.646	1	1.9	m	
EMAP Virginian Province	1990	VA90-134	15-AUG-1990	39.246	-76.557	1	9.2	m	
EMAP Virginian Province	1990	VA90-134	23-AUG-1990	39.246	-76.557	2	6.3	m	
EMAP Virginian Province	1990	VA90-134	06-SEP-1990	39.246	-76.557	3			
EMAP Virginian Province	1990	VA90-135	15-AUG-1990	39.219	-76.543	1			
EMAP Virginian Province	1990	VA90-136	05-AUG-1990	39.305	-76.41	1	3.4	m	
EMAP Virginian Province	1990	VA90-136	05-SEP-1990	39.305	-76.41	2			
EMAP Virginian Province	1990	VA90-137	05-AUG-1990	39.31	-76.409	1	3.6	m	
EMAP Virginian Province	1990	VA90-139	26-JUL-1990	39.255	-76.444	1			
EMAP Virginian Province	1990	VA90-140	15-AUG-1990	39.275	-76.45	1	1.8	m	
EMAP Virginian Province	1990	VA90-141	24-JUL-1990	37.675	-76.911	1	3.6	m	
EMAP Virginian Province	1990	VA90-141	04-SEP-1990	37.675	-76.911	2	4.0	m	
EMAP Virginian Province	1990	VA90-142	24-JUL-1990	37.528	-76.786	1	2.4	m	
EMAP Virginian Province	1990	VA90-143	24-JUL-1990	37.615	-76.847	1	9.8	m	
EMAP Virginian Province	1990	VA90-144	21-JUL-1990	37.13	-75.915	1	6.4	m	
EMAP Virginian Province	1990	VA90-145	21-JUL-1990	37.167	-75.921	1	1.5	m	
EMAP Virginian Province	1990	VA90-147	01-AUG-1990	40.75	-74.083	1	5.3	m	
EMAP Virginian Province	1990	VA90-150	19-JUL-1990	38.593	-75.112	1	1.7	m	
EMAP Virginian Province	1990	VA90-150	30-JUL-1990	38.593	-75.112	2	1.9	m	
EMAP Virginian Province	1990	VA90-150	08-AUG-1990	38.593	-75.112	3	1.8	m	
EMAP Virginian Province	1990	VA90-150	18-AUG-1990	38.593	-75.112	4	2.1	m	
EMAP Virginian Province	1990	VA90-150	28-AUG-1990	38.593	-75.112	5	1.9	m	
EMAP Virginian Province	1990	VA90-150	14-SEP-1990	38.593	-75.112	6	2.1	m	
EMAP Virginian Province	1990	VA90-151	19-JUL-1990	38.602	-75.129	1			
EMAP Virginian Province	1990	VA90-152	30-JUL-1990	38.584	-75.177	1	1.8	m	
EMAP Virginian Province	1990	VA90-153	30-JUL-1990	38.602	-75.137	1	2.7	m	
EMAP Virginian Province	1990	VA90-154	18-AUG-1990	38.595	-75.083	1	1.8	m	
EMAP Virginian Province	1990	VA90-155	30-JUL-1990	38.611	-75.11	1	2.0	m	
EMAP Virginian Province	1990	VA90-156	30-JUL-1990	41.0	-72.412	1	9.1	m	
EMAP Virginian Province	1990	VA90-156	09-SEP-1990	41.0	-72.412	2	9.9	m	
EMAP Virginian Province	1990	VA90-157	30-JUL-1990	41.0	-72.417	1	9.0	m	
EMAP Virginian Province	1990	VA90-158	10-AUG-1990	40.19	-74.032	1	2.9	m	
EMAP Virginian Province	1990	VA90-158	22-SEP-1990	40.19	-74.032	2			
EMAP Virginian Province	1990	VA90-159	19-JUL-1990	41.062	-72.002	1	16.4	m	
EMAP Virginian Province	1990	VA90-159	11-SEP-1990	41.062	-72.002	2	16.2	m	
EMAP Virginian Province	1990	VA90-160	19-JUL-1990	41.07	-72.035	1	15.3	m	
EMAP Virginian Province	1990	VA90-161	20-JUL-1990	40.872	-72.473	1	2.3	m	
EMAP Virginian Province	1990	VA90-161	10-SEP-1990	40.872	-72.473	2	3.1	m	
EMAP Virginian Province	1990	VA90-162	20-JUL-1990	40.86	-72.481	1	1.9	m	
EMAP Virginian Province	1990	VA90-164	01-AUG-1990	36.925	-76.345	1			
EMAP Virginian Province	1990	VA90-165	02-AUG-1990	36.852	-76.357	1	1.7	m	
EMAP Virginian Province	1990	VA90-166	27-JUL-1990	41.427	-70.517	1	9.0	m	
EMAP Virginian Province	1990	VA90-166	05-SEP-1990	41.427	-70.517	2	9.3	m	
EMAP Virginian Province	1990	VA90-167	27-JUL-1990	41.408	-70.482	1	10.0	m	
EMAP Virginian Province	1990	VA90-168	10-AUG-1990	40.193	-74.04	1			
EMAP Virginian Province	1990	VA90-169	21-AUG-1990	41.287	-73.072	1	6.0	m	
EMAP Virginian Province	1990	VA90-169	18-SEP-1990	41.287	-73.072	2	8.9	m	
EMAP Virginian Province	1990	VA90-170	21-AUG-1990	41.167	-73.092	1	6.7	m	
EMAP Virginian Province	1990	VA90-172	26-AUG-1990	38.859	-77.017	1	5.1	m	
EMAP Virginian Province	1990	VA90-173	30-JUL-1990	40.647	-74.058	1	13.6	m	
EMAP Virginian Province	1990	VA90-173	19-SEP-1990	40.647	-74.058	2	15.3	m	
EMAP Virginian Province	1990	VA90-174	20-JUL-1990	40.667	-74.045	1			
EMAP Virginian Province	1990	VA90-174	30-JUL-1990	40.667	-74.045	2	15.0	m	
EMAP Virginian Province	1990	VA90-177	12-AUG-1990	40.883	-73.943	1	3.6	m	
EMAP Virginian Province	1990	VA90-177	21-SEP-1990	40.883	-73.943	2	4.1	m	
EMAP Virginian Province	1990	VA90-178	19-AUG-1990	40.167	-74.728	1	6.6	m	
EMAP Virginian Province	1990	VA90-178	10-SEP-1990	40.167	-74.728	2	7.3	m	
EMAP Virginian Province	1990	VA90-179	19-AUG-1990	40.167	-74.729	1	3.8	m	
EMAP Virginian Province	1990	VA90-180	16-AUG-1990	38.07	-76.465	1	17.8	m	
EMAP Virginian Province	1990	VA90-180	15-SEP-1990	38.07	-76.465	2	17.1	m	
EMAP Virginian Province	1990	VA90-181	16-AUG-1990	38.051	-76.464	1			
EMAP Virginian Province	1990	VA90-182	06-AUG-1990	38.218	-76.786	1	10.2	m	
EMAP Virginian Province	1990	VA90-182	15-SEP-1990	38.218	-76.786	2	7.2	m	
EMAP Virginian Province	1990	VA90-183	06-AUG-1990	38.204	-76.786	1			
EMAP Virginian Province	1990	VA90-184	27-JUL-1990	38.398	-77.084	1	10.7	m	
EMAP Virginian Province	1990	VA90-184	06-AUG-1990	38.398	-77.084	2	9.1	m	
EMAP Virginian Province	1990	VA90-184	16-AUG-1990	38.398	-77.084	3	8.2	m	
EMAP Virginian Province	1990	VA90-184	25-AUG-1990	38.398	-77.084	4	6.7	m	
EMAP Virginian Province	1990	VA90-184	14-SEP-1990	38.398	-77.084	5			
EMAP Virginian Province	1990	VA90-185	27-JUL-1990	38.4	-77.083	1			
EMAP Virginian Province	1990	VA90-186	25-AUG-1990	38.5	-77.275	1	7.5	m	
EMAP Virginian Province	1990	VA90-186	14-SEP-1990	38.5	-77.275	2			
EMAP Virginian Province	1990	VA90-187	25-AUG-1990	38.5	-77.285	1	6.6	m	
EMAP Virginian Province	1990	VA90-188	26-AUG-1990	38.737	-77.033	1	9.7	m	
EMAP Virginian Province	1990	VA90-188	21-SEP-1990	38.737	-77.033	2	10.2	m	
EMAP Virginian Province	1990	VA90-189	26-AUG-1990	38.75	-77.036	1	2.3	m	
EMAP Virginian Province	1990	VA90-190	15-AUG-1990	37.737	-76.584	1	13.7	m	
EMAP Virginian Province	1990	VA90-190	07-SEP-1990	37.737	-76.584	2	15.9	m	
EMAP Virginian Province	1990	VA90-191	15-AUG-1990	37.733	-76.585	1	16.7	m	
EMAP Virginian Province	1990	VA90-192	26-JUL-1990	37.965	-76.867	1	2.4	m	
EMAP Virginian Province	1990	VA90-192	05-AUG-1990	37.965	-76.867	2	2.5	m	
EMAP Virginian Province	1990	VA90-192	15-AUG-1990	37.965	-76.867	3	2.4	m	
EMAP Virginian Province	1990	VA90-192	23-AUG-1990	37.965	-76.867	4	2.7	m	
EMAP Virginian Province	1990	VA90-192	07-SEP-1990	37.965	-76.867	5	2.5	m	
EMAP Virginian Province	1990	VA90-193	26-JUL-1990	37.967	-76.862	1	5.9	m	
EMAP Virginian Province	1990	VA90-194	26-JUL-1990	38.11	-77.0	1	8.5	m	
EMAP Virginian Province	1990	VA90-194	08-SEP-1990	38.11	-77.0	2	13.9	m	
EMAP Virginian Province	1990	VA90-195	26-JUL-1990	38.11	-77.0	1	14.2	m	
EMAP Virginian Province	1990	VA90-196	05-AUG-1990	38.165	-77.142	1	4.0	m	
EMAP Virginian Province	1990	VA90-196	08-SEP-1990	38.165	-77.142	2			
EMAP Virginian Province	1990	VA90-197	05-AUG-1990	38.167	-77.138	1	6.0	m	
EMAP Virginian Province	1990	VA90-198	12-AUG-1990	40.883	-73.933	1	8.3	m	
EMAP Virginian Province	1990	VA90-199	11-AUG-1990	41.15	-73.883	1	3.8	m	
EMAP Virginian Province	1990	VA90-199	20-SEP-1990	41.15	-73.883	2	2.3	m	
EMAP Virginian Province	1990	VA90-200	05-AUG-1990	38.2	-77.252	1	5.8	m	
EMAP Virginian Province	1990	VA90-200	08-SEP-1990	38.2	-77.252	2	4.9	m	
EMAP Virginian Province	1990	VA90-201	05-AUG-1990	38.2	-77.252	1	6.1	m	
EMAP Virginian Province	1990	VA90-202	02-AUG-1990	36.922	-76.351	1			
EMAP Virginian Province	1990	VA90-202	11-SEP-1990	36.922	-76.351	2	3.6	m	
EMAP Virginian Province	1990	VA90-203	01-AUG-1990	36.935	-76.351	1			
EMAP Virginian Province	1990	VA90-204	21-AUG-1990	37.032	-76.572	1	3.2	m	
EMAP Virginian Province	1990	VA90-204	10-SEP-1990	37.032	-76.572	2	2.8	m	
EMAP Virginian Province	1990	VA90-205	21-AUG-1990	37.033	-76.583	1	2.6	m	
EMAP Virginian Province	1990	VA90-206	22-AUG-1990	37.209	-76.798	1			
EMAP Virginian Province	1990	VA90-206	10-SEP-1990	37.209	-76.798	2	2.0	m	
EMAP Virginian Province	1990	VA90-207	22-AUG-1990	37.209	-76.792	1	2.4	m	
EMAP Virginian Province	1990	VA90-208	22-AUG-1990	37.27	-77.071	1			
EMAP Virginian Province	1990	VA90-208	10-SEP-1990	37.27	-77.071	2	9.9	m	
EMAP Virginian Province	1990	VA90-209	22-AUG-1990	37.268	-77.071	1	2.6	m	
EMAP Virginian Province	1990	VA90-210	23-JUL-1990	37.333	-77.273	1	4.1	m	
EMAP Virginian Province	1990	VA90-210	09-SEP-1990	37.333	-77.273	2	4.2	m	
EMAP Virginian Province	1990	VA90-212	11-AUG-1990	41.15	-73.896	1	10.7	m	
EMAP Virginian Province	1990	VA90-214	11-AUG-1990	41.383	-73.953	1	18.4	m	
EMAP Virginian Province	1990	VA90-215	10-AUG-1990	41.733	-73.945	1	15.2	m	
EMAP Virginian Province	1990	VA90-215	20-SEP-1990	41.733	-73.945	2	15.5	m	
EMAP Virginian Province	1990	VA90-216	10-AUG-1990	41.733	-73.943	1	14.4	m	
EMAP Virginian Province	1990	VA90-217	09-AUG-1990	42.0	-73.939	1	9.1	m	
EMAP Virginian Province	1990	VA90-217	19-SEP-1990	42.0	-73.939	2	8.3	m	
EMAP Virginian Province	1990	VA90-218	09-AUG-1990	42.0	-73.942	1	9.1	m	
EMAP Virginian Province	1990	VA90-219	28-JUL-1990	39.583	-75.582	1	3.1	m	
EMAP Virginian Province	1990	VA90-219	16-SEP-1990	39.583	-75.582	2	4.2	m	
EMAP Virginian Province	1990	VA90-220	18-AUG-1990	39.667	-75.535	1	12.0	m	
EMAP Virginian Province	1990	VA90-221	28-JUL-1990	39.583	-75.558	1	14.5	m	
EMAP Virginian Province	1990	VA90-221	26-AUG-1990	39.583	-75.558	2	13.0	m	
EMAP Virginian Province	1990	VA90-223	19-JUL-1990	39.75	-75.483	1	4.3	m	
EMAP Virginian Province	1990	VA90-223	29-JUL-1990	39.75	-75.483	2	4.6	m	
EMAP Virginian Province	1990	VA90-223	08-AUG-1990	39.75	-75.483	3	4.0	m	
EMAP Virginian Province	1990	VA90-223	18-AUG-1990	39.75	-75.483	4	4.0	m	
EMAP Virginian Province	1990	VA90-223	27-AUG-1990	39.75	-75.483	5	6.1	m	
EMAP Virginian Province	1990	VA90-223	11-SEP-1990	39.75	-75.483	6	5.2	m	
EMAP Virginian Province	1990	VA90-224	18-AUG-1990	39.847	-75.333	1	11.5	m	
EMAP Virginian Province	1990	VA90-225	29-JUL-1990	39.75	-75.488	1	12.0	m	
EMAP Virginian Province	1990	VA90-227	08-AUG-1990	39.881	-75.183	1	11.6	m	
EMAP Virginian Province	1990	VA90-227	11-SEP-1990	39.881	-75.183	2	14.4	m	
EMAP Virginian Province	1990	VA90-228	20-AUG-1990	39.974	-75.1	1	11.5	m	
EMAP Virginian Province	1990	VA90-229	08-AUG-1990	39.882	-75.183	1	13.6	m	
EMAP Virginian Province	1990	VA90-231	19-JUL-1990	40.05	-74.967	1	4.7	m	
EMAP Virginian Province	1990	VA90-231	10-SEP-1990	40.05	-74.967	2	5.2	m	
EMAP Virginian Province	1990	VA90-232	20-AUG-1990	40.1	-74.839	1	5.2	m	
EMAP Virginian Province	1990	VA90-233	19-JUL-1990	40.053	-74.967	1			
EMAP Virginian Province	1990	VA90-250	30-AUG-1990	39.277	-74.978	1			
EMAP Virginian Province	1990	VA90-250	09-SEP-1990	39.277	-74.978	2	8.0	m	
EMAP Virginian Province	1990	VA90-251	30-AUG-1990	39.212	-75.039	1			
EMAP Virginian Province	1990	VA90-252	26-AUG-1990	39.58	-75.495	1	4.1	m	
EMAP Virginian Province	1990	VA90-252	16-SEP-1990	39.58	-75.495	2	5.6	m	
EMAP Virginian Province	1990	VA90-253	26-AUG-1990	39.57	-75.514	1	5.8	m	
EMAP Virginian Province	1990	VA90-254	25-JUL-1990	39.48	-75.942	1	5.1	m	
EMAP Virginian Province	1990	VA90-254	15-SEP-1990	39.48	-75.942	3	4.1	m	
EMAP Virginian Province	1990	VA90-255	25-JUL-1990	39.428	-76.014	1	12.2	m	
EMAP Virginian Province	1990	VA90-256	22-JUL-1990	39.943	-74.102	1	1.8	m	
EMAP Virginian Province	1990	VA90-256	02-AUG-1990	39.943	-74.102	2	2.0	m	
EMAP Virginian Province	1990	VA90-256	10-AUG-1990	39.943	-74.102	3	1.9	m	
EMAP Virginian Province	1990	VA90-256	21-AUG-1990	39.943	-74.102	4	1.7	m	
EMAP Virginian Province	1990	VA90-256	27-AUG-1990	39.943	-74.102	5	2.0	m	
EMAP Virginian Province	1990	VA90-256	23-SEP-1990	39.943	-74.102	6			
EMAP Virginian Province	1990	VA90-257	22-JUL-1990	39.779	-74.125	1	3.5	m	
EMAP Virginian Province	1990	VA90-258	10-AUG-1990	37.3	-75.833	1	13.3	m	
EMAP Virginian Province	1990	VA90-259	10-AUG-1990	37.303	-75.802	1	5.8	m	
EMAP Virginian Province	1990	VA90-260	20-SEP-1990	40.705	-74.116	1	4.1	m	
EMAP Virginian Province	1991	VA91-025	06-AUG-1991	41.012	-73.242	1			
EMAP Virginian Province	1991	VA91-025	17-AUG-1991	41.012	-73.242	2	34.9	m	
EMAP Virginian Province	1991	VA91-025	18-AUG-1991	41.012	-73.242	3	31.0	m	
EMAP Virginian Province	1991	VA91-045	12-JUL-1991	38.161	-76.026	1	1.8	m	
EMAP Virginian Province	1991	VA91-045	15-JUL-1991	38.161	-76.026	2	2.0	m	
EMAP Virginian Province	1991	VA91-050	11-JUL-1991	38.012	-76.11	1	11.0	m	
EMAP Virginian Province	1991	VA91-050	12-JUL-1991	38.012	-76.11	2	10.8	m	
EMAP Virginian Province	1991	VA91-058	17-JUL-1991	39.129	-76.281	1	2.2	m	
EMAP Virginian Province	1991	VA91-058	18-JUL-1991	39.129	-76.281	2	2.1	m	
EMAP Virginian Province	1991	VA91-060	08-JUL-1991	37.715	-76.277	1	6.8	m	
EMAP Virginian Province	1991	VA91-060	09-JUL-1991	37.715	-76.277	2	6.7	m	
EMAP Virginian Province	1991	VA91-060	10-JUL-1991	37.715	-76.277	3	6.8	m	
EMAP Virginian Province	1991	VA91-079	05-AUG-1991	41.175	-72.706	1	30.0	m	
EMAP Virginian Province	1991	VA91-079	23-AUG-1991	41.175	-72.706	2	29.0	m	
EMAP Virginian Province	1991	VA91-079	25-AUG-1991	41.175	-72.706	3	30.0	m	
EMAP Virginian Province	1991	VA91-090	29-JUL-1991	39.27	-76.443	1	1.9	m	
EMAP Virginian Province	1991	VA91-090	31-JUL-1991	39.27	-76.443	2	1.7	m	
EMAP Virginian Province	1991	VA91-090	05-SEP-1991	39.27	-76.443	3	1.8	m	
EMAP Virginian Province	1991	VA91-136	29-JUL-1991	39.305	-76.41	1	3.2	m	
EMAP Virginian Province	1991	VA91-136	01-AUG-1991	39.305	-76.41	2	3.5	m	
EMAP Virginian Province	1991	VA91-150	22-AUG-1991	38.593	-75.112	1	2.0	m	
EMAP Virginian Province	1991	VA91-150	25-AUG-1991	38.593	-75.112	2	2.3	m	
EMAP Virginian Province	1991	VA91-173	03-AUG-1991	40.647	-74.058	1	15.0	m	
EMAP Virginian Province	1991	VA91-173	06-AUG-1991	40.647	-74.058	2	14.3	m	
EMAP Virginian Province	1991	VA91-188	22-JUL-1991	38.737	-77.033	1	5.0	m	
EMAP Virginian Province	1991	VA91-188	25-JUL-1991	38.737	-77.033	2	4.9	m	
EMAP Virginian Province	1991	VA91-215	28-AUG-1991	41.733	-73.945	1	16.2	m	
EMAP Virginian Province	1991	VA91-215	30-AUG-1991	41.733	-73.945	2	17.0	m	
EMAP Virginian Province	1991	VA91-261	03-AUG-1991	36.94	-76.214	1	5.4	m	
EMAP Virginian Province	1991	VA91-261	06-AUG-1991	36.94	-76.214	2	5.2	m	
EMAP Virginian Province	1991	VA91-262	15-AUG-1991	36.956	-76.008	1	21.8	m	
EMAP Virginian Province	1991	VA91-262	18-AUG-1991	36.956	-76.008	2	21.7	m	
EMAP Virginian Province	1991	VA91-263	03-AUG-1991	36.977	-76.483	1	3.5	m	
EMAP Virginian Province	1991	VA91-263	06-AUG-1991	36.977	-76.483	2	3.2	m	
EMAP Virginian Province	1991	VA91-265	15-AUG-1991	37.089	-76.132	1	12.9	m	
EMAP Virginian Province	1991	VA91-265	18-AUG-1991	37.089	-76.132	2	12.6	m	
EMAP Virginian Province	1991	VA91-266	17-AUG-1991	37.098	-76.333	1	2.2	m	
EMAP Virginian Province	1991	VA91-266	20-AUG-1991	37.098	-76.333	2	2.3	m	
EMAP Virginian Province	1991	VA91-267	17-AUG-1991	37.111	-76.297	1	5.6	m	
EMAP Virginian Province	1991	VA91-269	04-AUG-1991	37.163	-76.629	1	5.4	m	
EMAP Virginian Province	1991	VA91-269	07-AUG-1991	37.163	-76.629	2	5.5	m	
EMAP Virginian Province	1991	VA91-270	17-AUG-1991	37.221	-76.255	1	6.1	m	
EMAP Virginian Province	1991	VA91-270	20-AUG-1991	37.221	-76.255	2	6.6	m	
EMAP Virginian Province	1991	VA91-271	16-AUG-1991	37.237	-76.049	1	4.1	m	
EMAP Virginian Province	1991	VA91-271	19-AUG-1991	37.237	-76.049	2	4.7	m	
EMAP Virginian Province	1991	VA91-273	04-AUG-1991	37.241	-76.955	1	6.0	m	
EMAP Virginian Province	1991	VA91-273	07-AUG-1991	37.241	-76.955	2	6.6	m	
EMAP Virginian Province	1991	VA91-275	05-AUG-1991	37.32	-77.192	1	9.0	m	
EMAP Virginian Province	1991	VA91-275	08-AUG-1991	37.32	-77.192	2	7.4	m	
EMAP Virginian Province	1991	VA91-276	16-AUG-1991	37.37	-76.173	1	10.1	m	
EMAP Virginian Province	1991	VA91-276	20-AUG-1991	37.37	-76.173	2	10.7	m	
EMAP Virginian Province	1991	VA91-278	05-AUG-1991	37.379	-77.316	1	8.0	m	
EMAP Virginian Province	1991	VA91-278	08-AUG-1991	37.379	-77.316	2	8.1	m	
EMAP Virginian Province	1991	VA91-279	23-AUG-1991	37.518	-76.09	1	11.7	m	
EMAP Virginian Province	1991	VA91-279	26-AUG-1991	37.518	-76.09	2	11.6	m	
EMAP Virginian Province	1991	VA91-280	09-AUG-1991	37.533	-76.31	1	7.1	m	
EMAP Virginian Province	1991	VA91-281	09-AUG-1991	37.54	-76.405	1	5.7	m	
EMAP Virginian Province	1991	VA91-281	13-AUG-1991	37.54	-76.405	2	6.0	m	
EMAP Virginian Province	1991	VA91-282	09-AUG-1991	37.651	-76.215	1	11.4	m	
EMAP Virginian Province	1991	VA91-282	12-AUG-1991	37.651	-76.215	2	11.3	m	
EMAP Virginian Province	1991	VA91-283	23-AUG-1991	37.667	-76.007	1	14.9	m	
EMAP Virginian Province	1991	VA91-283	26-AUG-1991	37.667	-76.007	2	15.6	m	
EMAP Virginian Province	1991	VA91-284	10-AUG-1991	37.799	-76.131	1	10.3	m	
EMAP Virginian Province	1991	VA91-284	12-AUG-1991	37.799	-76.131	2	10.2	m	
EMAP Virginian Province	1991	VA91-285	22-AUG-1991	37.815	-75.924	1	4.8	m	
EMAP Virginian Province	1991	VA91-285	25-AUG-1991	37.815	-75.924	2	5.0	m	
EMAP Virginian Province	1991	VA91-286	11-AUG-1991	37.82	-76.298	1	7.1	m	
EMAP Virginian Province	1991	VA91-288	10-AUG-1991	37.831	-76.747	1	3.0	m	
EMAP Virginian Province	1991	VA91-288	13-AUG-1991	37.831	-76.747	2	3.0	m	
EMAP Virginian Province	1991	VA91-290	11-AUG-1991	37.85	-76.361	1	4.8	m	
EMAP Virginian Province	1991	VA91-290	13-AUG-1991	37.85	-76.361	2	4.5	m	
EMAP Virginian Province	1991	VA91-291	11-AUG-1991	37.931	-76.256	1	7.7	m	
EMAP Virginian Province	1991	VA91-291	13-AUG-1991	37.931	-76.256	2	7.6	m	
EMAP Virginian Province	1991	VA91-292	22-AUG-1991	37.947	-76.048	1	3.2	m	
EMAP Virginian Province	1991	VA91-292	25-AUG-1991	37.947	-76.048	2	4.2	m	
EMAP Virginian Province	1991	VA91-294	30-JUL-1991	38.039	-76.917	1	3.9	m	
EMAP Virginian Province	1991	VA91-294	02-AUG-1991	38.039	-76.917	2	3.9	m	
EMAP Virginian Province	1991	VA91-295	21-AUG-1991	38.08	-76.172	1	5.9	m	
EMAP Virginian Province	1991	VA91-295	24-AUG-1991	38.08	-76.172	2	6.1	m	
EMAP Virginian Province	1991	VA91-296	21-AUG-1991	38.096	-75.964	1	8.9	m	
EMAP Virginian Province	1991	VA91-296	24-AUG-1991	38.096	-75.964	2	8.9	m	
EMAP Virginian Province	1991	VA91-298	30-JUL-1991	38.14	-77.054	1	3.8	m	
EMAP Virginian Province	1991	VA91-298	02-AUG-1991	38.14	-77.054	2	4.1	m	
EMAP Virginian Province	1991	VA91-300	29-JUL-1991	38.181	-77.193	1	3.7	m	
EMAP Virginian Province	1991	VA91-300	01-AUG-1991	38.181	-77.193	2	4.5	m	
EMAP Virginian Province	1991	VA91-302	28-JUL-1991	38.207	-76.599	1	6.3	m	
EMAP Virginian Province	1991	VA91-302	31-JUL-1991	38.207	-76.599	2	6.3	m	
EMAP Virginian Province	1991	VA91-303	27-AUG-1991	38.212	-76.297	1	12.1	m	
EMAP Virginian Province	1991	VA91-303	28-AUG-1991	38.212	-76.297	2	12.2	m	
EMAP Virginian Province	1991	VA91-304	24-JUL-1991	38.222	-76.73	1	5.5	m	
EMAP Virginian Province	1991	VA91-305	23-AUG-1991	38.223	-75.217	1	1.9	m	
EMAP Virginian Province	1991	VA91-305	26-AUG-1991	38.223	-75.217	2	1.8	m	
EMAP Virginian Province	1991	VA91-306	28-JUL-1991	38.228	-76.697	1	5.4	m	
EMAP Virginian Province	1991	VA91-307	27-AUG-1991	38.228	-76.088	1	4.2	m	
EMAP Virginian Province	1991	VA91-307	28-AUG-1991	38.228	-76.088	2	4.1	m	
EMAP Virginian Province	1991	VA91-307	29-AUG-1991	38.228	-76.088	3	3.6	m	
EMAP Virginian Province	1991	VA91-308	29-AUG-1991	38.234	-75.992	1	5.1	m	
EMAP Virginian Province	1991	VA91-309	29-JUL-1991	38.235	-77.23	1	8.8	m	
EMAP Virginian Province	1991	VA91-309	01-AUG-1991	38.235	-77.23	2	7.9	m	
EMAP Virginian Province	1991	VA91-311	27-AUG-1991	38.249	-76.114	1	14.8	m	
EMAP Virginian Province	1991	VA91-311	28-AUG-1991	38.249	-76.114	2	8.8	m	
EMAP Virginian Province	1991	VA91-312	28-JUL-1991	38.256	-76.661	1	4.6	m	
EMAP Virginian Province	1991	VA91-314	24-JUL-1991	38.281	-76.711	1	2.2	m	
EMAP Virginian Province	1991	VA91-314	27-JUL-1991	38.281	-76.711	2	2.8	m	
EMAP Virginian Province	1991	VA91-315	24-JUL-1991	38.285	-76.928	1	3.3	m	
EMAP Virginian Province	1991	VA91-315	27-JUL-1991	38.285	-76.928	2	3.3	m	
EMAP Virginian Province	1991	VA91-316	27-AUG-1991	38.304	-76.184	1	2.8	m	
EMAP Virginian Province	1991	VA91-316	28-AUG-1991	38.304	-76.184	2	2.4	m	
EMAP Virginian Province	1991	VA91-316	29-AUG-1991	38.304	-76.184	3	2.6	m	
EMAP Virginian Province	1991	VA91-316	12-SEP-1991	38.304	-76.184	4	2.9	m	
EMAP Virginian Province	1991	VA91-317	29-AUG-1991	38.315	-76.02	1	3.9	m	
EMAP Virginian Province	1991	VA91-317	30-AUG-1991	38.315	-76.02	2	4.0	m	
EMAP Virginian Province	1991	VA91-318	23-AUG-1991	38.227	-75.177	1	1.8	m	
EMAP Virginian Province	1991	VA91-319	23-JUL-1991	38.336	-77.239	1	3.3	m	
EMAP Virginian Province	1991	VA91-319	26-JUL-1991	38.336	-77.239	2	3.3	m	
EMAP Virginian Province	1991	VA91-322	15-AUG-1991	38.519	-76.269	1	4.5	m	
EMAP Virginian Province	1991	VA91-322	18-AUG-1991	38.519	-76.269	2	5.0	m	
EMAP Virginian Province	1991	VA91-323	15-AUG-1991	38.549	-76.313	1	8.0	m	
EMAP Virginian Province	1991	VA91-325	15-AUG-1991	38.625	-76.464	1	11.2	m	
EMAP Virginian Province	1991	VA91-325	18-AUG-1991	38.625	-76.464	2	11.1	m	
EMAP Virginian Province	1991	VA91-326	23-JUL-1991	38.625	-77.162	1	3.9	m	
EMAP Virginian Province	1991	VA91-326	26-JUL-1991	38.625	-77.162	2	4.1	m	
EMAP Virginian Province	1991	VA91-327	24-AUG-1991	38.659	-75.097	1	2.2	m	
EMAP Virginian Province	1991	VA91-328	22-AUG-1991	38.675	-75.118	1	1.5	m	
EMAP Virginian Province	1991	VA91-328	24-AUG-1991	38.675	-75.118	2	1.7	m	
EMAP Virginian Province	1991	VA91-328	25-AUG-1991	38.675	-75.118	3	1.7	m	
EMAP Virginian Province	1991	VA91-330	17-AUG-1991	38.774	-76.185	1	9.4	m	
EMAP Virginian Province	1991	VA91-330	19-AUG-1991	38.774	-76.185	2	5.5	m	
EMAP Virginian Province	1991	VA91-331	16-AUG-1991	38.823	-76.218	1	10.1	m	
EMAP Virginian Province	1991	VA91-331	17-AUG-1991	38.823	-76.218	2	9.0	m	
EMAP Virginian Province	1991	VA91-332	16-AUG-1991	38.848	-76.203	1	12.0	m	
EMAP Virginian Province	1991	VA91-333	22-JUL-1991	38.859	-77.034	1	3.1	m	
EMAP Virginian Province	1991	VA91-333	25-JUL-1991	38.859	-77.034	2	3.8	m	
EMAP Virginian Province	1991	VA91-335	04-SEP-1991	38.864	-75.114	1	22.0	m	
EMAP Virginian Province	1991	VA91-335	06-SEP-1991	38.864	-75.114	2	24.0	m	
EMAP Virginian Province	1991	VA91-336	16-AUG-1991	38.906	-76.171	1	4.5	m	
EMAP Virginian Province	1991	VA91-336	19-AUG-1991	38.906	-76.171	2	4.3	m	
EMAP Virginian Province	1991	VA91-337	04-SEP-1991	38.997	-75.238	1	11.0	m	
EMAP Virginian Province	1991	VA91-337	06-SEP-1991	38.997	-75.238	2	10.8	m	
EMAP Virginian Province	1991	VA91-338	23-JUL-1991	39.011	-75.026	1	5.6	m	
EMAP Virginian Province	1991	VA91-338	26-JUL-1991	39.011	-75.026	2	6.2	m	
EMAP Virginian Province	1991	VA91-338	05-SEP-1991	39.011	-75.026	3	5.1	m	
EMAP Virginian Province	1991	VA91-339	28-JUL-1991	39.054	-76.421	1	4.0	m	
EMAP Virginian Province	1991	VA91-339	31-JUL-1991	39.054	-76.421	2	5.3	m	
EMAP Virginian Province	1991	VA91-340	04-SEP-1991	39.131	-75.362	1	4.4	m	
EMAP Virginian Province	1991	VA91-340	07-SEP-1991	39.131	-75.362	2	4.7	m	
EMAP Virginian Province	1991	VA91-341	22-JUL-1991	39.145	-75.15	1	3.5	m	
EMAP Virginian Province	1991	VA91-341	26-JUL-1991	39.145	-75.15	2	4.2	m	
EMAP Virginian Province	1991	VA91-341	05-SEP-1991	39.145	-75.15	3	4.5	m	
EMAP Virginian Province	1991	VA91-342	23-JUL-1991	39.158	-74.938	1	2.6	m	
EMAP Virginian Province	1991	VA91-342	26-JUL-1991	39.158	-74.938	2	2.6	m	
EMAP Virginian Province	1991	VA91-342	05-SEP-1991	39.158	-74.938	3	2.7	m	
EMAP Virginian Province	1991	VA91-343	28-JUL-1991	39.203	-76.336	1	5.0	m	
EMAP Virginian Province	1991	VA91-343	31-JUL-1991	39.203	-76.336	2	5.0	m	
EMAP Virginian Province	1991	VA91-343	05-SEP-1991	39.203	-76.336	3	4.9	m	
EMAP Virginian Province	1991	VA91-344	22-JUL-1991	39.278	-75.274	1	4.7	m	
EMAP Virginian Province	1991	VA91-344	26-JUL-1991	39.278	-75.274	2	6.2	m	
EMAP Virginian Province	1991	VA91-346	27-AUG-1991	39.37	-75.925	1	3.9	m	
EMAP Virginian Province	1991	VA91-346	29-AUG-1991	39.37	-75.925	2	3.8	m	
EMAP Virginian Province	1991	VA91-347	27-AUG-1991	39.38	-76.062	1	4.3	m	
EMAP Virginian Province	1991	VA91-348	24-JUL-1991	39.496	-74.382	1	1.6	m	
EMAP Virginian Province	1991	VA91-349	21-JUL-1991	39.504	-74.385	1	2.4	m	
EMAP Virginian Province	1991	VA91-349	24-JUL-1991	39.504	-74.385	2	2.1	m	
EMAP Virginian Province	1991	VA91-350	28-AUG-1991	39.533	-75.791	1	9.6	m	
EMAP Virginian Province	1991	VA91-351	30-JUL-1991	39.578	-76.091	1	9.9	m	
EMAP Virginian Province	1991	VA91-352	28-AUG-1991	39.555	-75.642	1	9.2	m	
EMAP Virginian Province	1991	VA91-352	30-AUG-1991	39.555	-75.642	2	11.2	m	
EMAP Virginian Province	1991	VA91-353	30-JUL-1991	39.588	-76.109	1	8.4	m	
EMAP Virginian Province	1991	VA91-353	01-AUG-1991	39.588	-76.109	2	9.3	m	
EMAP Virginian Province	1991	VA91-355	09-AUG-1991	39.667	-75.545	1	8.9	m	
EMAP Virginian Province	1991	VA91-355	12-AUG-1991	39.667	-75.545	2	8.7	m	
EMAP Virginian Province	1991	VA91-356	09-AUG-1991	39.717	-75.514	1	10.0	m	
EMAP Virginian Province	1991	VA91-357	09-AUG-1991	39.717	-75.572	1	4.2	m	
EMAP Virginian Province	1991	VA91-357	12-AUG-1991	39.717	-75.572	2	3.7	m	
EMAP Virginian Province	1991	VA91-358	10-AUG-1991	39.835	-75.351	1	3.9	m	
EMAP Virginian Province	1991	VA91-358	13-AUG-1991	39.835	-75.351	2	3.0	m	
EMAP Virginian Province	1991	VA91-360	10-AUG-1991	39.972	-75.1	1	11.5	m	
EMAP Virginian Province	1991	VA91-360	13-AUG-1991	39.972	-75.1	2	10.7	m	
EMAP Virginian Province	1991	VA91-362	05-AUG-1991	40.052	-74.111	1	2.5	m	
EMAP Virginian Province	1991	VA91-362	08-AUG-1991	40.052	-74.111	2	2.4	m	
EMAP Virginian Province	1991	VA91-363	05-AUG-1991	40.053	-74.067	1	1.8	m	
EMAP Virginian Province	1991	VA91-365	11-AUG-1991	40.101	-74.836	1	2.4	m	
EMAP Virginian Province	1991	VA91-365	13-AUG-1991	40.101	-74.836	2	2.7	m	
EMAP Virginian Province	1991	VA91-368	04-AUG-1991	40.49	-74.264	1	5.5	m	
EMAP Virginian Province	1991	VA91-369	04-AUG-1991	40.511	-74.3	1	7.5	m	
EMAP Virginian Province	1991	VA91-369	07-AUG-1991	40.511	-74.3	2	8.2	m	
EMAP Virginian Province	1991	VA91-370	04-AUG-1991	40.617	-73.888	1	5.6	m	
EMAP Virginian Province	1991	VA91-371	03-AUG-1991	40.616	-73.888	1	10.9	m	
EMAP Virginian Province	1991	VA91-371	07-AUG-1991	40.616	-73.888	2	11.1	m	
EMAP Virginian Province	1991	VA91-372	03-AUG-1991	40.642	-74.133	1	9.6	m	
EMAP Virginian Province	1991	VA91-372	06-AUG-1991	40.642	-74.133	2	10.7	m	
EMAP Virginian Province	1991	VA91-373	03-AUG-1991	40.648	-74.075	1	7.5	m	
EMAP Virginian Province	1991	VA91-375	05-AUG-1991	40.777	-73.855	1	5.7	m	
EMAP Virginian Province	1991	VA91-375	07-AUG-1991	40.777	-73.855	2	4.1	m	
EMAP Virginian Province	1991	VA91-376	06-AUG-1991	40.783	-73.939	1	6.6	m	
EMAP Virginian Province	1991	VA91-377	07-AUG-1991	40.792	-73.862	1	8.5	m	
EMAP Virginian Province	1991	VA91-378	04-AUG-1991	40.792	-73.932	1	8.3	m	
EMAP Virginian Province	1991	VA91-378	06-AUG-1991	40.792	-73.932	2	4.0	m	
EMAP Virginian Province	1991	VA91-379	05-AUG-1991	40.926	-73.619	1	15.1	m	
EMAP Virginian Province	1991	VA91-379	06-AUG-1991	40.926	-73.619	2	14.7	m	
EMAP Virginian Province	1991	VA91-380	17-AUG-1991	40.946	-73.181	1	14.6	m	
EMAP Virginian Province	1991	VA91-380	18-AUG-1991	40.946	-73.181	2	16.4	m	
EMAP Virginian Province	1991	VA91-381	15-AUG-1991	40.985	-72.419	1	16.7	m	
EMAP Virginian Province	1991	VA91-382	15-AUG-1991	41.0	-72.383	1	9.0	m	
EMAP Virginian Province	1991	VA91-384	27-AUG-1991	41.019	-73.893	1	5.9	m	
EMAP Virginian Province	1991	VA91-384	30-AUG-1991	41.019	-73.893	2	5.2	m	
EMAP Virginian Province	1991	VA91-385	22-AUG-1991	41.081	-73.304	1	15.5	m	
EMAP Virginian Province	1991	VA91-385	24-AUG-1991	41.081	-73.304	2	15.5	m	
EMAP Virginian Province	1991	VA91-386	06-AUG-1991	41.091	-73.084	1	37.0	m	
EMAP Virginian Province	1991	VA91-386	22-AUG-1991	41.091	-73.084	2	19.0	m	
EMAP Virginian Province	1991	VA91-386	24-AUG-1991	41.091	-73.084	3	33.0	m	
EMAP Virginian Province	1991	VA91-387	05-AUG-1991	41.1	-72.865	1	30.0	m	
EMAP Virginian Province	1991	VA91-387	23-AUG-1991	41.1	-72.865	2	30.0	m	
EMAP Virginian Province	1991	VA91-387	25-AUG-1991	41.1	-72.865	3	30.0	m	
EMAP Virginian Province	1991	VA91-388	05-AUG-1991	41.108	-72.645	1	30.0	m	
EMAP Virginian Province	1991	VA91-388	16-AUG-1991	41.108	-72.645	2	26.4	m	
EMAP Virginian Province	1991	VA91-388	18-AUG-1991	41.108	-72.645	3	26.3	m	
EMAP Virginian Province	1991	VA91-389	16-AUG-1991	41.116	-72.425	1	16.5	m	
EMAP Virginian Province	1991	VA91-389	18-AUG-1991	41.116	-72.425	2	17.5	m	
EMAP Virginian Province	1991	VA91-390	05-SEP-1991	41.131	-71.986	1	22.0	m	
EMAP Virginian Province	1991	VA91-390	07-SEP-1991	41.131	-71.986	2	21.0	m	
EMAP Virginian Province	1991	VA91-391	03-SEP-1991	41.138	-71.766	1	23.0	m	
EMAP Virginian Province	1991	VA91-391	05-SEP-1991	41.138	-71.766	2	24.0	m	
EMAP Virginian Province	1991	VA91-392	23-AUG-1991	41.244	-72.767	1	9.0	m	
EMAP Virginian Province	1991	VA91-392	25-AUG-1991	41.244	-72.767	2	8.0	m	
EMAP Virginian Province	1991	VA91-394	05-SEP-1991	41.268	-72.106	1	26.0	m	
EMAP Virginian Province	1991	VA91-394	07-SEP-1991	41.268	-72.106	2	24.0	m	
EMAP Virginian Province	1991	VA91-395	21-AUG-1991	41.283	-72.368	1	2.5	m	
EMAP Virginian Province	1991	VA91-397	27-AUG-1991	41.274	-73.967	1	8.7	m	
EMAP Virginian Province	1991	VA91-397	30-AUG-1991	41.274	-73.967	2	8.3	m	
EMAP Virginian Province	1991	VA91-398	11-AUG-1991	41.275	-71.886	1	43.0	m	
EMAP Virginian Province	1991	VA91-398	06-SEP-1991	41.275	-71.886	2	45.0	m	
EMAP Virginian Province	1991	VA91-398	08-SEP-1991	41.275	-71.886	3	40.0	m	
EMAP Virginian Province	1991	VA91-399	11-AUG-1991	41.282	-71.665	1	40.0	m	
EMAP Virginian Province	1991	VA91-399	06-SEP-1991	41.282	-71.665	2	40.0	m	
EMAP Virginian Province	1991	VA91-399	08-SEP-1991	41.282	-71.665	3	39.0	m	
EMAP Virginian Province	1991	VA91-400	25-JUL-1991	41.297	-70.099	1	6.5	m	
EMAP Virginian Province	1991	VA91-400	12-SEP-1991	41.297	-70.099	2	7.0	m	
EMAP Virginian Province	1991	VA91-401	04-SEP-1991	41.298	-72.183	1	9.5	m	
EMAP Virginian Province	1991	VA91-402	22-JUL-1991	41.316	-70.118	1	8.0	m	
EMAP Virginian Province	1991	VA91-402	23-JUL-1991	41.316	-70.118	2	8.0	m	
EMAP Virginian Province	1991	VA91-402	12-SEP-1991	41.316	-70.118	3	8.0	m	
EMAP Virginian Province	1991	VA91-403	21-AUG-1991	41.328	-72.353	1	4.0	m	
EMAP Virginian Province	1991	VA91-403	25-AUG-1991	41.328	-72.353	2	3.0	m	
EMAP Virginian Province	1991	VA91-404	22-JUL-1991	41.333	-70.017	1	6.0	m	
EMAP Virginian Province	1991	VA91-404	24-JUL-1991	41.333	-70.017	2	6.0	m	
EMAP Virginian Province	1991	VA91-405	04-SEP-1991	41.343	-72.179	1	3.1	m	
EMAP Virginian Province	1991	VA91-405	07-SEP-1991	41.343	-72.179	2	2.5	m	
EMAP Virginian Province	1991	VA91-406	29-JUL-1991	41.442	-70.9	1	14.0	m	
EMAP Virginian Province	1991	VA91-406	31-JUL-1991	41.442	-70.9	2	14.0	m	
EMAP Virginian Province	1991	VA91-407	29-JUL-1991	41.446	-70.679	1	9.0	m	
EMAP Virginian Province	1991	VA91-407	31-JUL-1991	41.446	-70.679	2	9.0	m	
EMAP Virginian Province	1991	VA91-408	30-JUL-1991	41.45	-70.457	1	8.0	m	
EMAP Virginian Province	1991	VA91-408	01-AUG-1991	41.45	-70.457	2	9.0	m	
EMAP Virginian Province	1991	VA91-409	22-JUL-1991	41.454	-70.235	1	14.1	m	
EMAP Virginian Province	1991	VA91-409	26-JUL-1991	41.454	-70.235	2	13.7	m	
EMAP Virginian Province	1991	VA91-410	09-AUG-1991	41.523	-71.065	1	5.0	m	
EMAP Virginian Province	1991	VA91-410	13-AUG-1991	41.523	-71.065	2	5.5	m	
EMAP Virginian Province	1991	VA91-411	28-AUG-1991	41.516	-73.992	1	9.0	m	
EMAP Virginian Province	1991	VA91-411	30-AUG-1991	41.516	-73.992	2	10.0	m	
EMAP Virginian Province	1991	VA91-413	09-AUG-1991	41.53	-71.094	1	3.0	m	
EMAP Virginian Province	1991	VA91-413	13-AUG-1991	41.53	-71.094	2	3.5	m	
EMAP Virginian Province	1991	VA91-414	28-JUL-1991	41.584	-70.797	1	12.0	m	
EMAP Virginian Province	1991	VA91-414	31-JUL-1991	41.584	-70.797	2	12.0	m	
EMAP Virginian Province	1991	VA91-414	13-SEP-1991	41.584	-70.797	3	13.0	m	
EMAP Virginian Province	1991	VA91-415	30-JUL-1991	41.592	-70.353	1	7.0	m	
EMAP Virginian Province	1991	VA91-415	01-AUG-1991	41.592	-70.353	2	7.0	m	
EMAP Virginian Province	1991	VA91-416	22-JUL-1991	41.596	-70.13	1	10.1	m	
EMAP Virginian Province	1991	VA91-416	26-JUL-1991	41.596	-70.13	2	9.6	m	
EMAP Virginian Province	1991	VA91-417	11-AUG-1991	41.641	-71.216	1	16.0	m	
EMAP Virginian Province	1991	VA91-418	11-AUG-1991	41.698	-71.206	1	6.5	m	
EMAP Virginian Province	1991	VA91-418	13-AUG-1991	41.698	-71.206	2	5.5	m	
EMAP Virginian Province	1991	VA91-419	10-AUG-1991	41.711	-71.164	1	6.5	m	
EMAP Virginian Province	1991	VA91-419	12-AUG-1991	41.711	-71.164	2	8.0	m	
EMAP Virginian Province	1991	VA91-421	10-AUG-1991	41.767	-71.123	1	7.5	m	
EMAP Virginian Province	1991	VA91-421	12-AUG-1991	41.767	-71.123	2	7.5	m	
EMAP Virginian Province	1991	VA91-422	29-AUG-1991	41.872	-73.935	1	13.1	m	
EMAP Virginian Province	1991	VA91-422	31-AUG-1991	41.872	-73.935	2	13.2	m	
EMAP Virginian Province	1991	VA91-424	29-AUG-1991	42.133	-73.907	1	6.8	m	
EMAP Virginian Province	1991	VA91-424	31-AUG-1991	42.133	-73.907	2	7.0	m	
EMAP Virginian Province	1991	VA91-426	10-JUL-1991	37.713	-76.275	1	9.6	m	
EMAP Virginian Province	1991	VA91-427	10-JUL-1991	37.709	-76.272	1	5.2	m	
EMAP Virginian Province	1991	VA91-428	10-JUL-1991	37.703	-76.267	1	6.2	m	
EMAP Virginian Province	1991	VA91-429	11-JUL-1991	38.006	-76.119	1	11.9	m	
EMAP Virginian Province	1991	VA91-430	11-JUL-1991	38.009	-76.115	1	11.6	m	
EMAP Virginian Province	1991	VA91-431	11-JUL-1991	38.0	-76.126	1	10.5	m	
EMAP Virginian Province	1991	VA91-432	16-JUL-1991	38.148	-76.012	1	2.6	m	
EMAP Virginian Province	1991	VA91-433	16-JUL-1991	38.151	-76.015	1	2.6	m	
EMAP Virginian Province	1991	VA91-434	16-JUL-1991	38.142	-76.007	1	2.6	m	
EMAP Virginian Province	1991	VA91-435	18-JUL-1991	39.124	-76.288	1	3.2	m	
EMAP Virginian Province	1991	VA91-436	17-JUL-1991	39.127	-76.284	1	3.3	m	
EMAP Virginian Province	1991	VA91-437	18-JUL-1991	39.12	-76.294	1	6.3	m	
EMAP Virginian Province	1992	VA92-025	04-AUG-1992	41.012	-73.242	1	34.8	m	
EMAP Virginian Province	1992	VA92-025	06-AUG-1992	41.012	-73.242	2	30.0	m	
EMAP Virginian Province	1992	VA92-025	26-AUG-1992	41.012	-73.242	1	36.5	m	
EMAP Virginian Province	1992	VA92-025	27-AUG-1992	41.012	-73.242	2	38.0	m	
EMAP Virginian Province	1992	VA92-045	02-AUG-1992	38.161	-76.026	1	1.7	m	
EMAP Virginian Province	1992	VA92-045	27-AUG-1992	38.161	-76.026	2	1.9	m	
EMAP Virginian Province	1992	VA92-050	03-AUG-1992	38.012	-76.11	1	10.7	m	
EMAP Virginian Province	1992	VA92-050	27-AUG-1992	38.012	-76.11	2	9.8	m	
EMAP Virginian Province	1992	VA92-058	03-AUG-1992	39.129	-76.281	1	2.3	m	
EMAP Virginian Province	1992	VA92-058	30-AUG-1992	39.129	-76.281	2	2.0	m	
EMAP Virginian Province	1992	VA92-060	05-AUG-1992	37.715	-76.277	1	6.4	m	
EMAP Virginian Province	1992	VA92-060	30-AUG-1992	37.715	-76.277	2	6.8	m	
EMAP Virginian Province	1992	VA92-079	10-AUG-1992	41.175	-72.706	1	27.3	m	
EMAP Virginian Province	1992	VA92-079	11-AUG-1992	41.175	-72.706	2	28.0	m	
EMAP Virginian Province	1992	VA92-079	26-AUG-1992	41.175	-72.706	3	28.0	m	
EMAP Virginian Province	1992	VA92-079	09-SEP-1992	41.175	-72.706	4	28.0	m	
EMAP Virginian Province	1992	VA92-136	04-AUG-1992	39.305	-76.41	1	2.8	m	
EMAP Virginian Province	1992	VA92-136	29-AUG-1992	39.305	-76.41	2	3.8	m	
EMAP Virginian Province	1992	VA92-150	17-AUG-1992	38.593	-75.112	1	1.7	m	
EMAP Virginian Province	1992	VA92-150	27-AUG-1992	38.593	-75.112	2	2.0	m	
EMAP Virginian Province	1992	VA92-173	27-JUL-1992	40.647	-74.058	1	15.1	m	
EMAP Virginian Province	1992	VA92-173	24-AUG-1992	40.647	-74.058	2	15.0	m	
EMAP Virginian Province	1992	VA92-178	31-JUL-1992	40.167	-74.728	1	6.6	m	
EMAP Virginian Province	1992	VA92-178	23-AUG-1992	40.167	-74.728	2	5.1	m	
EMAP Virginian Province	1992	VA92-188	27-JUL-1992	38.737	-77.033	1	5.7	m	
EMAP Virginian Province	1992	VA92-188	26-AUG-1992	38.737	-77.033	2	5.1	m	
EMAP Virginian Province	1992	VA92-215	12-AUG-1992	41.733	-73.945	1	16.7	m	
EMAP Virginian Province	1992	VA92-215	23-AUG-1992	41.733	-73.945	2	15.9	m	
EMAP Virginian Province	1992	VA92-451	10-AUG-1992	36.864	-76.519	1	2.5	m	
EMAP Virginian Province	1992	VA92-452	09-AUG-1992	36.881	-76.012	1	3.2	m	
EMAP Virginian Province	1992	VA92-453	10-AUG-1992	36.927	-76.417	1	5.0	m	
EMAP Virginian Province	1992	VA92-454	08-AUG-1992	37.015	-76.173	1	6.3	m	
EMAP Virginian Province	1992	VA92-455	08-AUG-1992	37.031	-75.967	1	5.6	m	
EMAP Virginian Province	1992	VA92-456	15-AUG-1992	37.057	-76.62	1	3.1	m	
EMAP Virginian Province	1992	VA92-457	15-AUG-1992	37.087	-76.599	1	4.0	m	
EMAP Virginian Province	1992	VA92-460	11-AUG-1992	37.163	-76.091	1	8.6	m	
EMAP Virginian Province	1992	VA92-461	14-AUG-1992	37.226	-76.895	1	4.1	m	
EMAP Virginian Province	1992	VA92-462	11-AUG-1992	37.295	-76.214	1	10.0	m	
EMAP Virginian Province	1992	VA92-464	17-AUG-1992	37.312	-77.106	1	7.7	m	
EMAP Virginian Province	1992	VA92-465	21-AUG-1992	37.329	-76.381	1	5.7	m	
EMAP Virginian Province	1992	VA92-466	21-AUG-1992	37.331	-76.394	1	5.7	m	
EMAP Virginian Province	1992	VA92-467	16-AUG-1992	37.318	-77.284	1	2.7	m	
EMAP Virginian Province	1992	VA92-468	14-AUG-1992	37.345	-76.874	1	5.1	m	
EMAP Virginian Province	1992	VA92-469	16-AUG-1992	37.356	-77.271	1	6.1	m	
EMAP Virginian Province	1992	VA92-470	23-AUG-1992	37.444	-76.132	1	11.7	m	
EMAP Virginian Province	1992	VA92-471	18-AUG-1992	37.561	-76.905	1	5.0	m	
EMAP Virginian Province	1992	VA92-472	23-AUG-1992	37.576	-76.256	1	7.4	m	
EMAP Virginian Province	1992	VA92-473	22-AUG-1992	37.592	-76.049	1	14.7	m	
EMAP Virginian Province	1992	VA92-474	22-AUG-1992	37.725	-76.173	1	16.6	m	
EMAP Virginian Province	1992	VA92-475	24-AUG-1992	37.741	-75.966	1	6.8	m	
EMAP Virginian Province	1992	VA92-476	04-AUG-1992	37.807	-76.682	1	3.1	m	
EMAP Virginian Province	1992	VA92-477	04-AUG-1992	37.811	-76.694	1	4.3	m	
EMAP Virginian Province	1992	VA92-478	24-AUG-1992	37.873	-76.09	1	10.7	m	
EMAP Virginian Province	1992	VA92-481	06-AUG-1992	37.984	-76.906	1	2.1	m	
EMAP Virginian Province	1992	VA92-482	30-AUG-1992	38.006	-76.214	1	21.6	m	
EMAP Virginian Province	1992	VA92-483	15-AUG-1992	38.064	-75.793	1	3.3	m	
EMAP Virginian Province	1992	VA92-484	06-AUG-1992	38.095	-77.035	1	6.8	m	
EMAP Virginian Province	1992	VA92-484	29-AUG-1992	38.095	-77.035	2	6.5	m	
EMAP Virginian Province	1992	VA92-485	28-AUG-1992	38.124	-76.498	1	5.5	m	
EMAP Virginian Province	1992	VA92-486	28-AUG-1992	38.134	-76.483	1	4.8	m	
EMAP Virginian Province	1992	VA92-486	31-AUG-1992	38.134	-76.483	2	4.3	m	
EMAP Virginian Province	1992	VA92-487	02-AUG-1992	38.154	-76.13	1	6.8	m	
EMAP Virginian Province	1992	VA92-488	15-AUG-1992	38.215	-75.851	1	2.7	m	
EMAP Virginian Province	1992	VA92-489	30-JUL-1992	38.213	-76.92	1	4.7	m	
EMAP Virginian Province	1992	VA92-490	30-JUL-1992	38.245	-76.811	1	2.0	m	
EMAP Virginian Province	1992	VA92-491	14-AUG-1992	38.286	-76.255	1	6.1	m	
EMAP Virginian Province	1992	VA92-492	31-JUL-1992	38.346	-76.854	1	3.0	m	
EMAP Virginian Province	1992	VA92-493	29-JUL-1992	38.354	-77.193	1	9.6	m	
EMAP Virginian Province	1992	VA92-494	29-JUL-1992	38.396	-77.325	1	3.3	m	
EMAP Virginian Province	1992	VA92-495	16-AUG-1992	38.402	-75.088	1	2.4	m	
EMAP Virginian Province	1992	VA92-496	16-AUG-1992	38.418	-75.093	1	2.0	m	
EMAP Virginian Province	1992	VA92-497	14-AUG-1992	38.419	-76.381	1	15.1	m	
EMAP Virginian Province	1992	VA92-499	28-JUL-1992	38.618	-77.212	1	2.7	m	
EMAP Virginian Province	1992	VA92-500	30-AUG-1992	38.699	-76.422	1	19.3	m	
EMAP Virginian Province	1992	VA92-501	28-AUG-1992	38.742	-76.31	1	2.4	m	
EMAP Virginian Province	1992	VA92-502	27-JUL-1992	38.778	-77.036	1	2.5	m	
EMAP Virginian Province	1992	VA92-503	18-AUG-1992	38.924	-75.282	1	2.4	m	
EMAP Virginian Province	1992	VA92-504	06-AUG-1992	38.922	-76.492	1	3.9	m	
EMAP Virginian Province	1992	VA92-505	10-AUG-1992	38.938	-75.07	1	13.4	m	
EMAP Virginian Province	1992	VA92-506	06-AUG-1992	38.98	-76.476	1	4.7	m	
EMAP Virginian Province	1992	VA92-507	02-AUG-1992	39.066	-76.44	1	4.0	m	
EMAP Virginian Province	1992	VA92-508	12-AUG-1992	39.071	-75.194	1	8.6	m	
EMAP Virginian Province	1992	VA92-509	09-AUG-1992	39.092	-74.767	1	1.3	m	
EMAP Virginian Province	1992	VA92-510	10-AUG-1992	39.085	-74.982	1	5.9	m	
EMAP Virginian Province	1992	VA92-511	03-AUG-1992	39.128	-76.379	1	5.8	m	
EMAP Virginian Province	1992	VA92-512	09-AUG-1992	39.18	-74.7	1	3.1	m	
EMAP Virginian Province	1992	VA92-513	26-AUG-1992	39.204	-75.318	1	7.0	m	
EMAP Virginian Province	1992	VA92-514	04-AUG-1992	39.277	-76.293	1	3.7	m	
EMAP Virginian Province	1992	VA92-515	08-AUG-1992	39.293	-74.613	1	4.3	m	
EMAP Virginian Province	1992	VA92-516	08-AUG-1992	39.323	-74.668	1	4.4	m	
EMAP Virginian Province	1992	VA92-517	26-AUG-1992	39.338	-75.443	1	9.0	m	
EMAP Virginian Province	1992	VA92-518	11-AUG-1992	39.382	-75.348	1	7.6	m	
EMAP Virginian Province	1992	VA92-519	05-AUG-1992	39.428	-76.24	1	1.7	m	
EMAP Virginian Province	1992	VA92-520	20-AUG-1992	39.471	-75.568	1	9.9	m	
EMAP Virginian Province	1992	VA92-521	28-AUG-1992	39.479	-75.897	1	2.2	m	
EMAP Virginian Province	1992	VA92-522	20-AUG-1992	39.642	-75.584	1	7.2	m	
EMAP Virginian Province	1992	VA92-523	21-AUG-1992	39.791	-75.43	1	5.5	m	
EMAP Virginian Province	1992	VA92-524	21-AUG-1992	39.816	-75.387	1	15.1	m	
EMAP Virginian Province	1992	VA92-525	22-AUG-1992	39.944	-75.135	1	14.2	m	
EMAP Virginian Province	1992	VA92-526	22-AUG-1992	40.072	-74.919	1	3.6	m	
EMAP Virginian Province	1992	VA92-527	30-JUL-1992	40.092	-74.079	1	2.0	m	
EMAP Virginian Province	1992	VA92-528	29-JUL-1992	40.495	-74.193	1	3.5	m	
EMAP Virginian Province	1992	VA92-529	29-JUL-1992	40.502	-74.191	1	5.0	m	
EMAP Virginian Province	1992	VA92-530	28-JUL-1992	40.693	-74.118	1	3.6	m	
EMAP Virginian Province	1992	VA92-532	27-AUG-1992	40.792	-72.718	1	1.9	m	
EMAP Virginian Province	1992	VA92-533	02-AUG-1992	40.83	-73.717	1	2.5	m	
EMAP Virginian Province	1992	VA92-534	02-AUG-1992	40.857	-73.667	1	7.0	m	
EMAP Virginian Province	1992	VA92-535	03-AUG-1992	40.91	-73.36	1	3.2	m	
EMAP Virginian Province	1992	VA92-536	03-AUG-1992	40.967	-73.105	1	7.9	m	
EMAP Virginian Province	1992	VA92-537	21-AUG-1992	40.979	-73.904	1	5.7	m	
EMAP Virginian Province	1992	VA92-538	20-AUG-1992	40.999	-73.571	1	6.0	m	
EMAP Virginian Province	1992	VA92-539	04-AUG-1992	41.009	-73.352	1	40.1	m	
EMAP Virginian Province	1992	VA92-539	07-AUG-1992	41.009	-73.352	2	40.0	m	
EMAP Virginian Province	1992	VA92-540	28-AUG-1992	41.02	-72.19	1	3.3	m	
EMAP Virginian Province	1992	VA92-541	06-AUG-1992	41.027	-72.914	1	39.3	m	
EMAP Virginian Province	1992	VA92-542	06-AUG-1992	41.018	-73.133	1	44.1	m	
EMAP Virginian Province	1992	VA92-542	07-AUG-1992	41.018	-73.133	2	48.0	m	
EMAP Virginian Province	1992	VA92-543	29-AUG-1992	41.039	-72.33	1	11.8	m	
EMAP Virginian Province	1992	VA92-544	08-AUG-1992	41.036	-72.694	1	29.1	m	
EMAP Virginian Province	1992	VA92-544	10-AUG-1992	41.036	-72.694	2	27.0	m	
EMAP Virginian Province	1992	VA92-545	28-AUG-1992	41.066	-71.921	1	2.0	m	
EMAP Virginian Province	1992	VA92-546	29-AUG-1992	41.091	-72.367	1	4.7	m	
EMAP Virginian Province	1992	VA92-547	11-AUG-1992	41.163	-73.036	1	13.4	m	
EMAP Virginian Province	1992	VA92-548	10-AUG-1992	41.181	-72.596	1	28.0	m	
EMAP Virginian Province	1992	VA92-549	08-AUG-1992	41.172	-72.816	1	18.8	m	
EMAP Virginian Province	1992	VA92-549	11-AUG-1992	41.172	-72.816	2	19.0	m	
EMAP Virginian Province	1992	VA92-550	17-AUG-1992	41.196	-72.156	1	23.8	m	
EMAP Virginian Province	1992	VA92-551	10-AUG-1992	41.189	-72.376	1	46.4	m	
EMAP Virginian Province	1992	VA92-552	21-AUG-1992	41.192	-73.956	1	1.8	m	
EMAP Virginian Province	1992	VA92-553	15-AUG-1992	41.21	-71.715	1	27.7	m	
EMAP Virginian Province	1992	VA92-553	18-AUG-1992	41.21	-71.715	2	33.0	m	
EMAP Virginian Province	1992	VA92-554	15-AUG-1992	41.203	-71.936	1	35.9	m	
EMAP Virginian Province	1992	VA92-554	18-AUG-1992	41.203	-71.936	2	30.3	m	
EMAP Virginian Province	1992	VA92-555	22-AUG-1992	41.235	-73.949	1	6.3	m	
EMAP Virginian Province	1992	VA92-556	14-AUG-1992	41.353	-71.685	1	1.5	m	
EMAP Virginian Province	1992	VA92-557	28-JUL-1992	41.383	-70.287	1	5.0	m	
EMAP Virginian Province	1992	VA92-558	28-JUL-1992	41.387	-70.066	1	12.4	m	
EMAP Virginian Province	1992	VA92-558	29-JUL-1992	41.387	-70.066	2	13.8	m	
EMAP Virginian Province	1992	VA92-559	14-AUG-1992	41.4	-71.506	1	2.0	m	
EMAP Virginian Province	1992	VA92-560	22-AUG-1992	41.472	-73.994	1	3.4	m	
EMAP Virginian Province	1992	VA92-561	16-AUG-1992	41.513	-70.85	1	17.0	m	
EMAP Virginian Province	1992	VA92-562	29-JUL-1992	41.525	-70.183	1	9.2	m	
EMAP Virginian Province	1992	VA92-563	31-JUL-1992	41.521	-70.405	1	12.1	m	
EMAP Virginian Province	1992	VA92-564	30-JUL-1992	41.517	-70.627	1	13.1	m	
EMAP Virginian Province	1992	VA92-565	30-JUL-1992	41.579	-70.522	1	2.3	m	
EMAP Virginian Province	1992	VA92-566	15-AUG-1992	41.583	-71.233	1	4.9	m	
EMAP Virginian Province	1992	VA92-567	31-JUL-1992	41.64	-70.258	1	3.2	m	
EMAP Virginian Province	1992	VA92-568	16-AUG-1992	41.655	-70.745	1	6.8	m	
EMAP Virginian Province	1992	VA92-569	27-JUL-1992	41.68	-69.941	1	4.7	m	
EMAP Virginian Province	1992	VA92-570	23-AUG-1992	41.801	-73.948	1	12.4	m	
EMAP Virginian Province	1992	VA92-571	24-AUG-1992	42.088	-73.929	1	11.6	m	
EMAP Virginian Province	1993	VA93-025	01-AUG-1993	41.012	-73.242	1	36.0	m	
EMAP Virginian Province	1993	VA93-025	31-AUG-1993	41.012	-73.242	2	35.0	m	
EMAP Virginian Province	1993	VA93-045	07-AUG-1993	38.161	-76.026	1	1.4	m	
EMAP Virginian Province	1993	VA93-045	01-SEP-1993	38.161	-76.026	2	2.0	m	
EMAP Virginian Province	1993	VA93-050	29-JUL-1993	38.012	-76.11	1	10.2	m	
EMAP Virginian Province	1993	VA93-050	26-AUG-1993	38.012	-76.11	2	11.0	m	
EMAP Virginian Province	1993	VA93-058	04-AUG-1993	39.129	-76.281	1	2.3	m	
EMAP Virginian Province	1993	VA93-058	02-SEP-1993	39.129	-76.281	2	2.2	m	
EMAP Virginian Province	1993	VA93-060	07-AUG-1993	37.715	-76.277	1	7.2	m	
EMAP Virginian Province	1993	VA93-060	26-AUG-1993	37.715	-76.277	2	6.2	m	
EMAP Virginian Province	1993	VA93-079	03-AUG-1993	41.175	-72.706	1	28.0	m	
EMAP Virginian Province	1993	VA93-079	01-SEP-1993	41.175	-72.706	2	28.0	m	
EMAP Virginian Province	1993	VA93-136	03-AUG-1993	39.305	-76.41	1	3.4	m	
EMAP Virginian Province	1993	VA93-136	30-AUG-1993	39.305	-76.41	2	3.6	m	
EMAP Virginian Province	1993	VA93-150	13-AUG-1993	38.593	-75.112	1	2.0	m	
EMAP Virginian Province	1993	VA93-150	02-SEP-1993	38.593	-75.112	2	1.0	m	
EMAP Virginian Province	1993	VA93-173	07-AUG-1993	40.647	-74.058	1	15.3	m	
EMAP Virginian Province	1993	VA93-173	02-SEP-1993	40.647	-74.058	2	15.8	m	
EMAP Virginian Province	1993	VA93-178	27-JUL-1993	40.167	-74.728	1	6.3	m	
EMAP Virginian Province	1993	VA93-178	31-AUG-1993	40.167	-74.728	2	3.8	m	
EMAP Virginian Province	1993	VA93-188	02-AUG-1993	38.737	-77.033	1	1.9	m	
EMAP Virginian Province	1993	VA93-188	25-AUG-1993	38.737	-77.033	2	5.2	m	
EMAP Virginian Province	1993	VA93-215	27-JUL-1993	41.733	-73.945	1	15.0	m	
EMAP Virginian Province	1993	VA93-215	28-JUL-1993	41.733	-73.945	2	12.5	m	
EMAP Virginian Province	1993	VA93-215	03-SEP-1993	41.733	-73.945	3	6.0	m	
EMAP Virginian Province	1993	VA93-601	18-SEP-1993	36.948	-76.111	1	9.0	m	
EMAP Virginian Province	1993	VA93-602	13-AUG-1993	37.007	-76.533	1	3.2	m	
EMAP Virginian Province	1993	VA93-604	26-JUL-1993	37.097	-76.029	1	4.3	m	
EMAP Virginian Province	1993	VA93-606	14-AUG-1993	37.201	-76.689	1	4.1	m	
EMAP Virginian Province	1993	VA93-607	27-AUG-1993	37.213	-76.358	1	5.8	m	
EMAP Virginian Province	1993	VA93-608	04-SEP-1993	37.229	-76.152	1	10.1	m	
EMAP Virginian Province	1993	VA93-609	15-AUG-1993	37.302	-77.0	1	12.1	m	
EMAP Virginian Province	1993	VA93-610	16-AUG-1993	37.307	-77.25	1	5.5	m	
EMAP Virginian Province	1993	VA93-611	28-AUG-1993	37.343	-76.624	1	4.4	m	
EMAP Virginian Province	1993	VA93-612	04-SEP-1993	37.378	-76.07	1	13.7	m	
EMAP Virginian Province	1993	VA93-613	17-AUG-1993	37.404	-77.394	1	9.0	m	
EMAP Virginian Province	1993	VA93-615	04-SEP-1993	37.51	-76.194	1	9.5	m	
EMAP Virginian Province	1993	VA93-616	27-JUL-1993	37.526	-75.987	1	6.2	m	
EMAP Virginian Province	1993	VA93-616	28-JUL-1993	37.526	-75.987	2	6.0	m	
EMAP Virginian Province	1993	VA93-617	22-AUG-1993	37.642	-76.318	1	4.3	m	
EMAP Virginian Province	1993	VA93-618	03-SEP-1993	37.659	-76.111	1	13.0	m	
EMAP Virginian Province	1993	VA93-619	28-JUL-1993	37.675	-75.904	1	3.0	m	
EMAP Virginian Province	1993	VA93-620	08-AUG-1993	37.708	-76.482	1	5.6	m	
EMAP Virginian Province	1993	VA93-621	20-AUG-1993	37.943	-76.846	1	2.3	m	
EMAP Virginian Province	1993	VA93-622	07-AUG-1993	37.791	-76.235	1	10.8	m	
EMAP Virginian Province	1993	VA93-623	08-AUG-1993	37.807	-76.028	1	4.7	m	
EMAP Virginian Province	1993	VA93-624	08-AUG-1993	37.823	-75.82	1	5.0	m	
EMAP Virginian Province	1993	VA93-626	03-SEP-1993	37.939	-76.152	1	19.0	m	
EMAP Virginian Province	1993	VA93-627	09-AUG-1993	37.955	-75.944	1	18.9	m	
EMAP Virginian Province	1993	VA93-628	19-AUG-1993	38.087	-76.982	1	4.5	m	
EMAP Virginian Province	1993	VA93-630	04-AUG-1993	38.072	-76.277	1	11.3	m	
EMAP Virginian Province	1993	VA93-631	09-AUG-1993	38.088	-76.068	1	3.1	m	
EMAP Virginian Province	1993	VA93-632	20-AUG-1993	38.162	-77.088	1	7.8	m	
EMAP Virginian Province	1993	VA93-633	01-SEP-1993	38.129	-75.89	1	2.9	m	
EMAP Virginian Province	1993	VA93-634	17-AUG-1993	38.148	-75.233	1	2.3	m	
EMAP Virginian Province	1993	VA93-635	23-AUG-1993	38.2	-77.223	1	5.5	m	
EMAP Virginian Province	1993	VA93-637	11-AUG-1993	38.22	-76.701	1	7.2	m	
EMAP Virginian Province	1993	VA93-638	30-JUL-1993	38.22	-76.193	1	6.1	m	
EMAP Virginian Province	1993	VA93-639	21-AUG-1993	38.249	-77.264	1	6.2	m	
EMAP Virginian Province	1993	VA93-640	10-AUG-1993	38.25	-75.842	1	2.3	m	
EMAP Virginian Province	1993	VA93-641	16-AUG-1993	38.317	-75.109	1	2.2	m	
EMAP Virginian Province	1993	VA93-642	10-AUG-1993	38.328	-75.895	1	2.1	m	
EMAP Virginian Province	1993	VA93-643	09-AUG-1993	38.344	-76.981	1	4.6	m	
EMAP Virginian Province	1993	VA93-644	02-SEP-1993	38.353	-76.318	1	39.0	m	
EMAP Virginian Province	1993	VA93-645	10-AUG-1993	38.419	-77.273	1	6.1	m	
EMAP Virginian Province	1993	VA93-647	05-AUG-1993	38.485	-76.444	1	11.5	m	
EMAP Virginian Province	1993	VA93-648	05-AUG-1993	38.486	-76.659	1	4.6	m	
EMAP Virginian Province	1993	VA93-649	27-AUG-1993	38.597	-76.065	1	3.8	m	
EMAP Virginian Province	1993	VA93-650	29-AUG-1993	38.633	-76.359	1	4.1	m	
EMAP Virginian Province	1993	VA93-651	01-AUG-1993	38.685	-77.104	1	1.6	m	
EMAP Virginian Province	1993	VA93-652	28-AUG-1993	38.715	-76.114	1	1.9	m	
EMAP Virginian Province	1993	VA93-653	27-AUG-1993	38.765	-76.485	1	8.9	m	
EMAP Virginian Province	1993	VA93-654	15-AUG-1993	38.857	-75.22	1	2.7	m	
EMAP Virginian Province	1993	VA93-655	03-AUG-1993	38.903	-77.073	1	4.6	m	
EMAP Virginian Province	1993	VA93-657	25-AUG-1993	38.914	-76.401	1	16.9	m	
EMAP Virginian Province	1993	VA93-658	26-AUG-1993	38.92	-76.28	1	5.8	m	
EMAP Virginian Province	1993	VA93-659	21-AUG-1993	38.95	-74.895	1	2.8	m	
EMAP Virginian Province	1993	VA93-660	22-AUG-1993	39.004	-75.132	1	4.4	m	
EMAP Virginian Province	1993	VA93-661	05-AUG-1993	39.025	-76.188	1	10.6	m	
EMAP Virginian Province	1993	VA93-663	19-AUG-1993	39.138	-75.256	1	6.2	m	
EMAP Virginian Province	1993	VA93-664	19-AUG-1993	39.152	-75.044	1	3.3	m	
EMAP Virginian Province	1993	VA93-666	14-AUG-1993	39.271	-75.381	1	6.0	m	
EMAP Virginian Province	1993	VA93-667	02-AUG-1993	39.359	-76.144	1	7.9	m	
EMAP Virginian Province	1993	VA93-668	30-JUL-1993	39.404	-75.506	1	12.0	m	
EMAP Virginian Province	1993	VA93-669	22-AUG-1993	39.407	-74.465	1	1.5	m	
EMAP Virginian Province	1993	VA93-670	01-AUG-1993	39.48	-76.07	1	3.8	m	
EMAP Virginian Province	1993	VA93-671	21-AUG-1993	39.558	-74.32	1	2.5	m	
EMAP Virginian Province	1993	VA93-672	01-AUG-1993	39.567	-75.959	1	2.5	m	
EMAP Virginian Province	1993	VA93-673	29-JUL-1993	39.712	-75.496	1	2.6	m	
EMAP Virginian Province	1993	VA93-675	28-JUL-1993	39.867	-75.214	1	14.4	m	
EMAP Virginian Province	1993	VA93-676	20-AUG-1993	39.945	-74.183	1	2.1	m	
EMAP Virginian Province	1993	VA93-677	26-JUL-1993	40.142	-74.733	1	2.9	m	
EMAP Virginian Province	1993	VA93-678	27-JUL-1993	40.018	-75.033	1	5.8	m	
EMAP Virginian Province	1993	VA93-681	09-AUG-1993	40.533	-74.073	1	4.6	m	
EMAP Virginian Province	1993	VA93-682	08-AUG-1993	40.55	-74.248	1	7.8	m	
EMAP Virginian Province	1993	VA93-683	11-AUG-1993	40.649	-73.476	1	2.7	m	
EMAP Virginian Province	1993	VA93-684	07-AUG-1993	40.74	-74.118	1	2.8	m	
EMAP Virginian Province	1993	VA93-685	10-AUG-1993	40.772	-73.759	1	2.0	m	
EMAP Virginian Province	1993	VA93-686	01-SEP-1993	40.898	-73.515	1	7.0	m	
EMAP Virginian Province	1993	VA93-687	31-AUG-1993	40.931	-73.509	1	14.0	m	
EMAP Virginian Province	1993	VA93-688	31-AUG-1993	40.941	-73.291	1	11.0	m	
EMAP Virginian Province	1993	VA93-689	28-AUG-1993	41.013	-72.048	1	2.2	m	
EMAP Virginian Province	1993	VA93-690	27-AUG-1993	41.059	-72.148	1	6.3	m	
EMAP Virginian Province	1993	VA93-693	30-JUL-1993	41.086	-73.194	1	18.7	m	
EMAP Virginian Province	1993	VA93-694	26-JUL-1993	41.088	-73.899	1	3.7	m	
EMAP Virginian Province	1993	VA93-695	02-AUG-1993	41.095	-72.975	1	26.0	m	
EMAP Virginian Province	1993	VA93-695	03-AUG-1993	41.095	-72.975	2	26.0	m	
EMAP Virginian Province	1993	VA93-696	02-AUG-1993	41.104	-72.755	1	30.0	m	
EMAP Virginian Province	1993	VA93-697	04-AUG-1993	41.113	-72.535	1	30.0	m	
EMAP Virginian Province	1993	VA93-698	27-AUG-1993	41.128	-72.096	1	12.2	m	
EMAP Virginian Province	1993	VA93-699	17-SEP-1993	41.135	-71.876	1	29.1	m	
EMAP Virginian Province	1993	VA93-700	17-SEP-1993	41.142	-71.655	1	21.0	m	
EMAP Virginian Province	1993	VA93-702	26-AUG-1993	41.246	-72.937	1	3.8	m	
EMAP Virginian Province	1993	VA93-703	25-AUG-1993	41.249	-72.657	1	8.1	m	
EMAP Virginian Province	1993	VA93-704	25-AUG-1993	41.257	-72.437	1	9.4	m	
EMAP Virginian Province	1993	VA93-705	05-AUG-1993	41.265	-72.216	1	30.0	m	
EMAP Virginian Province	1993	VA93-706	16-SEP-1993	41.279	-71.775	1	40.0	m	
EMAP Virginian Province	1993	VA93-707	17-SEP-1993	41.285	-71.555	1	42.4	m	
EMAP Virginian Province	1993	VA93-709	13-AUG-1993	41.327	-71.94	1	6.1	m	
EMAP Virginian Province	1993	VA93-710	26-JUL-1993	41.331	-73.977	1	27.3	m	
EMAP Virginian Province	1993	VA93-711	19-AUG-1993	41.336	-70.773	1	6.6	m	
EMAP Virginian Province	1993	VA93-712	14-AUG-1993	41.347	-71.715	1	2.8	m	
EMAP Virginian Province	1993	VA93-713	13-AUG-1993	41.351	-72.091	1	4.9	m	
EMAP Virginian Province	1993	VA93-714	19-AUG-1993	41.388	-70.463	1	3.4	m	
EMAP Virginian Province	1993	VA93-715	14-SEP-1993	41.444	-70.789	1	16.0	m	
EMAP Virginian Province	1993	VA93-716	14-SEP-1993	41.452	-70.346	1	16.0	m	
EMAP Virginian Province	1993	VA93-717	15-SEP-1993	41.456	-70.124	1	13.0	m	
EMAP Virginian Province	1993	VA93-718	14-AUG-1993	41.571	-71.351	1	10.5	m	
EMAP Virginian Province	1993	VA93-719	27-JUL-1993	41.578	-73.954	1	18.6	m	
EMAP Virginian Province	1993	VA93-720	16-AUG-1993	41.582	-70.908	1	6.5	m	
EMAP Virginian Province	1993	VA93-721	20-AUG-1993	41.586	-70.686	1	14.6	m	
EMAP Virginian Province	1993	VA93-722	21-AUG-1993	41.595	-70.465	1	2.0	m	
EMAP Virginian Province	1993	VA93-723	22-AUG-1993	41.594	-70.242	1	6.1	m	
EMAP Virginian Province	1993	VA93-724	22-AUG-1993	41.597	-70.019	1	5.9	m	
EMAP Virginian Province	1993	VA93-725	15-AUG-1993	41.812	-71.398	1	13.0	m	
EMAP Virginian Province	1993	VA93-726	28-JUL-1993	41.936	-73.948	1	6.5	m	
EMAP Virginian Province	1993	VA93-727	29-JUL-1993	42.192	-73.858	1	13.0	m	
EMAP Virginian Province	1993	VA93-728	15-AUG-1993	37.289	-76.992	1	4.2	m	
EMAP Virginian Province	1993	VA93-729	28-AUG-1993	37.525	-76.788	1	3.0	m	
EMAP Virginian Province	1993	VA93-730	08-AUG-1993	37.683	-76.464	1	5.3	m	
EMAP Virginian Province	1993	VA93-731	19-AUG-1993	38.081	-76.956	1	3.2	m	
EMAP Virginian Province	1993	VA93-732	17-AUG-1993	38.326	-75.1	1	3.4	m	
EMAP Virginian Province	1993	VA93-733	02-AUG-1993	38.901	-77.066	1	5.6	m	
EMAP Virginian Province	1993	VA93-734	26-JUL-1993	40.128	-74.742	1	2.0	m	
EMAP Virginian Province	1993	VA93-735	07-AUG-1993	40.647	-74.18	1	2.3	m	
EMAP Virginian Province	1993	VA93-735	08-AUG-1993	40.647	-74.18	2	3.8	m	
EMAP Virginian Province	1993	VA93-736	27-JUL-1993	41.557	-73.982	1	12.7	m	
EMAP Virginian Province	1993	VA93-737	15-AUG-1993	41.721	-71.363	1	3.1	m	
